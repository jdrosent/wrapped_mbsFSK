* NGSPICE file created from wrapped_mbsFSK.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

.subckt wrapped_mbsFSK active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12] la1_data_in[13] la1_data_in[14]
+ la1_data_in[15] la1_data_in[16] la1_data_in[17] la1_data_in[18] la1_data_in[19]
+ la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22] la1_data_in[23] la1_data_in[24]
+ la1_data_in[25] la1_data_in[26] la1_data_in[27] la1_data_in[28] la1_data_in[29]
+ la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3] la1_data_in[4] la1_data_in[5]
+ la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9] la1_data_out[0] la1_data_out[10]
+ la1_data_out[11] la1_data_out[12] la1_data_out[13] la1_data_out[14] la1_data_out[15]
+ la1_data_out[16] la1_data_out[17] la1_data_out[18] la1_data_out[19] la1_data_out[1]
+ la1_data_out[20] la1_data_out[21] la1_data_out[22] la1_data_out[23] la1_data_out[24]
+ la1_data_out[25] la1_data_out[26] la1_data_out[27] la1_data_out[28] la1_data_out[29]
+ la1_data_out[2] la1_data_out[30] la1_data_out[31] la1_data_out[3] la1_data_out[4]
+ la1_data_out[5] la1_data_out[6] la1_data_out[7] la1_data_out[8] la1_data_out[9]
+ la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12] la1_oenb[13] la1_oenb[14] la1_oenb[15]
+ la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19] la1_oenb[1] la1_oenb[20] la1_oenb[21]
+ la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25] la1_oenb[26] la1_oenb[27] la1_oenb[28]
+ la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31] la1_oenb[3] la1_oenb[4] la1_oenb[5]
+ la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9] vccd1 vssd1 wb_clk_i
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3155_ _3157_/CLK _3155_/D vssd1 vssd1 vccd1 vccd1 _3155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2106_ _1765_/X _2848_/B _1980_/C vssd1 vssd1 vccd1 vccd1 _2106_/Y sky130_fd_sc_hd__a21oi_1
X_3086_ _3086_/CLK _3086_/D vssd1 vssd1 vccd1 vccd1 _3086_/Q sky130_fd_sc_hd__dfxtp_1
X_2037_ _1795_/X _1953_/X _2223_/B vssd1 vssd1 vccd1 vccd1 _2547_/C sky130_fd_sc_hd__a21oi_2
XFILLER_22_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2939_ _3408_/A _2939_/B vssd1 vssd1 vccd1 vccd1 _2940_/A sky130_fd_sc_hd__and2_1
XFILLER_2_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_26 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_52 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_450 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_188 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_62 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2724_ _2471_/B _2471_/C _2471_/D _2275_/X vssd1 vssd1 vccd1 vccd1 _2724_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2655_ _2570_/X _2654_/Y _2649_/X vssd1 vssd1 vccd1 vccd1 _3163_/D sky130_fd_sc_hd__a21oi_1
X_1606_ _1606_/A vssd1 vssd1 vccd1 vccd1 _1611_/A sky130_fd_sc_hd__buf_4
X_2586_ _2783_/A vssd1 vssd1 vccd1 vccd1 _2586_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1537_ _1661_/A vssd1 vssd1 vccd1 vccd1 _1669_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3207_ _3230_/CLK _3207_/D vssd1 vssd1 vccd1 vccd1 _3207_/Q sky130_fd_sc_hd__dfxtp_1
X_3138_ _3268_/CLK _3138_/D vssd1 vssd1 vccd1 vccd1 _3138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3069_ _3069_/CLK _3069_/D vssd1 vssd1 vccd1 vccd1 _3069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_383 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2440_ _3109_/Q _2432_/X _2435_/X _3108_/Q vssd1 vssd1 vccd1 vccd1 _2440_/Y sky130_fd_sc_hd__a22oi_1
X_2371_ _3084_/Q _2365_/X _2368_/X _3083_/Q vssd1 vssd1 vccd1 vccd1 _2371_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_342 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2707_ _3178_/Q _2842_/B vssd1 vssd1 vccd1 vccd1 _2707_/X sky130_fd_sc_hd__or2_1
X_2638_ _2638_/A vssd1 vssd1 vccd1 vccd1 _2638_/X sky130_fd_sc_hd__clkbuf_2
X_2569_ _2567_/X _2568_/Y _2479_/X vssd1 vssd1 vccd1 vccd1 _3136_/D sky130_fd_sc_hd__a21oi_1
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_61 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_71 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1940_ _1940_/A vssd1 vssd1 vccd1 vccd1 _2046_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1871_ _2268_/A _1981_/A _1895_/A vssd1 vssd1 vccd1 vccd1 _2546_/C sky130_fd_sc_hd__a21oi_1
XFILLER_50_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2423_ _3102_/Q _2418_/X _2422_/X _3101_/Q vssd1 vssd1 vccd1 vccd1 _2423_/Y sky130_fd_sc_hd__a22oi_1
X_2354_ _2406_/A vssd1 vssd1 vccd1 vccd1 _2354_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2285_ _2283_/X _2284_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _3053_/D sky130_fd_sc_hd__o21a_1
XFILLER_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2070_ _2819_/A _2152_/A _2211_/B _2915_/B vssd1 vssd1 vccd1 vccd1 _2072_/A sky130_fd_sc_hd__or4_2
XFILLER_81_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2972_ _1696_/A _2987_/Q _2113_/A _2971_/X vssd1 vssd1 vccd1 vccd1 _3268_/D sky130_fd_sc_hd__o211a_1
X_1923_ _2178_/A _1843_/B _2268_/B vssd1 vssd1 vccd1 vccd1 _2170_/C sky130_fd_sc_hd__a21oi_2
X_1854_ _2801_/B _1852_/Y _1853_/X vssd1 vssd1 vccd1 vccd1 _2995_/D sky130_fd_sc_hd__a21oi_1
X_3365__7 vssd1 vssd1 vccd1 vccd1 _3365__7/HI _3365_/A sky130_fd_sc_hd__conb_1
X_1785_ _1777_/Y _1784_/Y _1672_/B vssd1 vssd1 vccd1 vccd1 _2992_/D sky130_fd_sc_hd__a21oi_1
X_3455_ _3455_/A _1629_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
X_2406_ _2406_/A vssd1 vssd1 vccd1 vccd1 _2406_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3386_ _3386_/A _1587_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
X_2337_ _2351_/A vssd1 vssd1 vccd1 vccd1 _2337_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2268_ _2268_/A _2268_/B vssd1 vssd1 vccd1 vccd1 _2269_/D sky130_fd_sc_hd__nor2_1
XFILLER_72_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2199_ _2686_/B _2199_/B vssd1 vssd1 vccd1 vccd1 _2500_/C sky130_fd_sc_hd__nand2_1
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3080_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1570_ _1574_/A vssd1 vssd1 vccd1 vccd1 _1570_/Y sky130_fd_sc_hd__inv_2
XANTENNA_5 _1661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_56 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3244_/CLK _3240_/D vssd1 vssd1 vccd1 vccd1 _3240_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3241_/CLK _3171_/D vssd1 vssd1 vccd1 vccd1 _3171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_404 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2122_ _2819_/A _2122_/B _2152_/A _2566_/B vssd1 vssd1 vccd1 vccd1 _2122_/X sky130_fd_sc_hd__or4b_1
XFILLER_66_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_278 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2053_ _2046_/A _2677_/B _2756_/A _2778_/B _2756_/C vssd1 vssd1 vccd1 vccd1 _2053_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_34_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2955_ _2960_/A _3261_/Q vssd1 vssd1 vccd1 vccd1 _2955_/X sky130_fd_sc_hd__or2_1
X_1906_ _3000_/Q _1863_/X _1874_/X _2999_/Q vssd1 vssd1 vccd1 vccd1 _1906_/Y sky130_fd_sc_hd__a22oi_1
X_2886_ _3232_/Q _2761_/X _2528_/X _3231_/Q _2524_/A vssd1 vssd1 vccd1 vccd1 _2886_/X
+ sky130_fd_sc_hd__o221a_1
X_1837_ _1893_/B _1960_/D _2034_/D _1960_/B vssd1 vssd1 vccd1 vccd1 _1887_/B sky130_fd_sc_hd__nand4b_4
X_1768_ _1890_/D _1953_/B vssd1 vssd1 vccd1 vccd1 _1951_/B sky130_fd_sc_hd__nand2_1
X_1699_ _2508_/A vssd1 vssd1 vccd1 vccd1 _2959_/A sky130_fd_sc_hd__clkbuf_2
X_3438_ _3438_/A _1611_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _3369_/A _1566_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2740_ _2769_/A _2740_/B _2740_/C vssd1 vssd1 vccd1 vccd1 _2741_/A sky130_fd_sc_hd__and3_1
X_2671_ _2761_/A vssd1 vssd1 vccd1 vccd1 _2671_/X sky130_fd_sc_hd__clkbuf_2
X_1622_ _1624_/A vssd1 vssd1 vccd1 vccd1 _1622_/Y sky130_fd_sc_hd__inv_2
X_1553_ _1556_/A vssd1 vssd1 vccd1 vccd1 _1553_/Y sky130_fd_sc_hd__inv_2
X_3223_ _3231_/CLK _3223_/D vssd1 vssd1 vccd1 vccd1 _3223_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3154_ _3154_/CLK _3154_/D vssd1 vssd1 vccd1 vccd1 _3154_/Q sky130_fd_sc_hd__dfxtp_1
X_2105_ _2105_/A _2105_/B vssd1 vssd1 vccd1 vccd1 _2105_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3085_ _3086_/CLK _3085_/D vssd1 vssd1 vccd1 vccd1 _3085_/Q sky130_fd_sc_hd__dfxtp_1
X_2036_ _2036_/A _2170_/D _1804_/X vssd1 vssd1 vccd1 vccd1 _2756_/C sky130_fd_sc_hd__or3b_2
X_3445__71 vssd1 vssd1 vccd1 vccd1 _3445__71/HI _3445_/A sky130_fd_sc_hd__conb_1
XFILLER_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2938_ _2938_/A vssd1 vssd1 vccd1 vccd1 _3254_/D sky130_fd_sc_hd__clkbuf_1
X_2869_ _3225_/Q _2853_/X _2859_/X _3224_/Q vssd1 vssd1 vccd1 vccd1 _2869_/Y sky130_fd_sc_hd__a22oi_1
X_3373__15 vssd1 vssd1 vccd1 vccd1 _3373__15/HI _3373_/A sky130_fd_sc_hd__conb_1
XFILLER_77_38 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2723_ _3182_/Q _2512_/X _2483_/X _3181_/Q _2722_/X vssd1 vssd1 vccd1 vccd1 _3182_/D
+ sky130_fd_sc_hd__o221a_1
X_2654_ _3163_/Q _2653_/X _2642_/X _3162_/Q vssd1 vssd1 vccd1 vccd1 _2654_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_8_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1605_ _1605_/A vssd1 vssd1 vccd1 vccd1 _1605_/Y sky130_fd_sc_hd__inv_2
X_2585_ _2585_/A vssd1 vssd1 vccd1 vccd1 _2783_/A sky130_fd_sc_hd__buf_2
X_1536_ input1/X vssd1 vssd1 vccd1 vccd1 _1661_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3206_ _3234_/CLK _3206_/D vssd1 vssd1 vccd1 vccd1 _3206_/Q sky130_fd_sc_hd__dfxtp_1
X_3137_ _3157_/CLK _3137_/D vssd1 vssd1 vccd1 vccd1 _3137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3068_ _3194_/CLK _3068_/D vssd1 vssd1 vccd1 vccd1 _3068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2019_ _2871_/A vssd1 vssd1 vccd1 vccd1 _2019_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_159 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2370_ _2131_/Y _2369_/Y _2362_/X vssd1 vssd1 vccd1 vccd1 _3083_/D sky130_fd_sc_hd__a21oi_1
XFILLER_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2706_ _2619_/D _2477_/D _2519_/D _3177_/Q _1705_/A vssd1 vssd1 vccd1 vccd1 _2706_/X
+ sky130_fd_sc_hd__o32a_1
X_2637_ _1899_/Y _2636_/Y _2621_/X vssd1 vssd1 vccd1 vccd1 _3157_/D sky130_fd_sc_hd__a21oi_1
X_2568_ _3136_/Q _2556_/X _2559_/X _3135_/Q vssd1 vssd1 vccd1 vccd1 _2568_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2499_ _1999_/A _2274_/B _2061_/X vssd1 vssd1 vccd1 vccd1 _2500_/D sky130_fd_sc_hd__a21oi_1
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1870_ _2178_/A vssd1 vssd1 vccd1 vccd1 _1981_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_450 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2422_ _2559_/A vssd1 vssd1 vccd1 vccd1 _2422_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2353_ _2166_/Y _2352_/Y _2349_/X vssd1 vssd1 vccd1 vccd1 _3077_/D sky130_fd_sc_hd__a21oi_1
XFILLER_69_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2284_ _3053_/Q _2081_/X _2020_/X _3052_/Q vssd1 vssd1 vccd1 vccd1 _2284_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_310 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1999_ _1999_/A _2274_/B vssd1 vssd1 vccd1 vccd1 _2778_/B sky130_fd_sc_hd__and2_1
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_54 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2971_ _2971_/A _3268_/Q vssd1 vssd1 vccd1 vccd1 _2971_/X sky130_fd_sc_hd__or2_1
X_1922_ _1965_/A vssd1 vssd1 vccd1 vccd1 _2268_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_42_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1853_ _2942_/A vssd1 vssd1 vccd1 vccd1 _1853_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1784_ _2992_/Q _2773_/A _1783_/X _2991_/Q vssd1 vssd1 vccd1 vccd1 _1784_/Y sky130_fd_sc_hd__a22oi_1
X_3454_ _3454_/A _1627_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
X_2405_ _2054_/Y _2404_/Y _2401_/X vssd1 vssd1 vccd1 vccd1 _3095_/D sky130_fd_sc_hd__a21oi_1
X_3385_ _3385_/A _1586_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2336_ _2201_/X _2334_/Y _2335_/X vssd1 vssd1 vccd1 vccd1 _3071_/D sky130_fd_sc_hd__a21oi_1
XFILLER_57_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2267_ _2267_/A _2267_/B vssd1 vssd1 vccd1 vccd1 _2819_/B sky130_fd_sc_hd__and2_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_90 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2198_ _2198_/A _2198_/B vssd1 vssd1 vccd1 vccd1 _2205_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3379__21 vssd1 vssd1 vccd1 vccd1 _3379__21/HI _3379_/A sky130_fd_sc_hd__conb_1
XFILLER_61_73 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _2471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_68 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3244_/CLK _3170_/D vssd1 vssd1 vccd1 vccd1 _3170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2121_ _2119_/X _2120_/Y _2092_/X vssd1 vssd1 vccd1 vccd1 _3023_/D sky130_fd_sc_hd__a21oi_1
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2052_ _2049_/X _2051_/Y _2043_/X vssd1 vssd1 vccd1 vccd1 _3012_/D sky130_fd_sc_hd__a21oi_1
XFILLER_22_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2954_ _2954_/A vssd1 vssd1 vccd1 vccd1 _2954_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_382 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1905_ _2157_/C _1904_/Y _1861_/X vssd1 vssd1 vccd1 vccd1 _1905_/Y sky130_fd_sc_hd__o21ai_2
X_2885_ _2885_/A _2885_/B _2885_/C vssd1 vssd1 vccd1 vccd1 _2885_/X sky130_fd_sc_hd__or3_1
X_1836_ _1836_/A vssd1 vssd1 vccd1 vccd1 _1893_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1767_ _1888_/B vssd1 vssd1 vccd1 vccd1 _1953_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1698_ _2550_/A vssd1 vssd1 vccd1 vccd1 _2508_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3437_ _3437_/A _1610_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3368_/A _1565_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2319_ _3065_/Q _2311_/X _2314_/X _3064_/Q vssd1 vssd1 vccd1 vccd1 _2319_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2670_ _2670_/A vssd1 vssd1 vccd1 vccd1 _3168_/D sky130_fd_sc_hd__clkbuf_1
X_1621_ _1624_/A vssd1 vssd1 vccd1 vccd1 _1621_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1552_ _1556_/A vssd1 vssd1 vccd1 vccd1 _1552_/Y sky130_fd_sc_hd__inv_2
X_3222_ _3232_/CLK _3222_/D vssd1 vssd1 vccd1 vccd1 _3222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3153_ _3157_/CLK _3153_/D vssd1 vssd1 vccd1 vccd1 _3153_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2104_ _2100_/Y _2103_/Y _2092_/X vssd1 vssd1 vccd1 vccd1 _3020_/D sky130_fd_sc_hd__a21oi_1
XFILLER_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3084_ _3086_/CLK _3084_/D vssd1 vssd1 vccd1 vccd1 _3084_/Q sky130_fd_sc_hd__dfxtp_1
X_2035_ _2061_/C _2035_/B _2034_/D vssd1 vssd1 vccd1 vccd1 _2170_/D sky130_fd_sc_hd__nor3b_2
XFILLER_35_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_102 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2937_ _3407_/A _2939_/B vssd1 vssd1 vccd1 vccd1 _2938_/A sky130_fd_sc_hd__and2_1
XFILLER_50_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3460__86 vssd1 vssd1 vccd1 vccd1 _3460__86/HI _3460_/A sky130_fd_sc_hd__conb_1
X_2868_ _2175_/X _2866_/Y _2867_/X vssd1 vssd1 vccd1 vccd1 _3224_/D sky130_fd_sc_hd__a21oi_1
X_1819_ _2477_/B vssd1 vssd1 vccd1 vccd1 _1819_/X sky130_fd_sc_hd__buf_2
X_2799_ _2929_/B vssd1 vssd1 vccd1 vccd1 _2907_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2722_ _2935_/B vssd1 vssd1 vccd1 vccd1 _2722_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2653_ _2829_/A vssd1 vssd1 vccd1 vccd1 _2653_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1604_ _1605_/A vssd1 vssd1 vccd1 vccd1 _1604_/Y sky130_fd_sc_hd__inv_2
X_2584_ _2584_/A _2584_/B _2693_/C _2584_/D vssd1 vssd1 vccd1 vccd1 _2584_/X sky130_fd_sc_hd__or4_4
X_3205_ _3230_/CLK _3205_/D vssd1 vssd1 vccd1 vccd1 _3205_/Q sky130_fd_sc_hd__dfxtp_1
X_3136_ _3157_/CLK _3136_/D vssd1 vssd1 vccd1 vccd1 _3136_/Q sky130_fd_sc_hd__dfxtp_1
X_3067_ _3070_/CLK _3067_/D vssd1 vssd1 vccd1 vccd1 _3067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2018_ _2848_/B _1831_/D _2015_/X _2017_/X vssd1 vssd1 vccd1 vccd1 _2018_/X sky130_fd_sc_hd__o31a_1
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3092_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3430__56 vssd1 vssd1 vccd1 vccd1 _3430__56/HI _3430_/A sky130_fd_sc_hd__conb_1
X_2705_ _2704_/B _2703_/X _2704_/Y _1681_/A vssd1 vssd1 vccd1 vccd1 _3177_/D sky130_fd_sc_hd__a211oi_1
X_2636_ _3157_/Q _2635_/X _2611_/X _3156_/Q vssd1 vssd1 vccd1 vccd1 _2636_/Y sky130_fd_sc_hd__a22oi_1
X_2567_ _2848_/A _2912_/A _2567_/C _2716_/B vssd1 vssd1 vccd1 vccd1 _2567_/X sky130_fd_sc_hd__or4_4
X_2498_ _2638_/A vssd1 vssd1 vccd1 vccd1 _2498_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3119_ _3154_/CLK _3119_/D vssd1 vssd1 vccd1 vccd1 _3119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3470_ _3470_/A _1650_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
X_2421_ _2585_/A vssd1 vssd1 vccd1 vccd1 _2559_/A sky130_fd_sc_hd__buf_2
X_2352_ _3077_/Q _2351_/X _2341_/X _3076_/Q vssd1 vssd1 vccd1 vccd1 _2352_/Y sky130_fd_sc_hd__a22oi_1
X_2283_ _2223_/Y _2780_/A _2181_/B _2017_/X vssd1 vssd1 vccd1 vccd1 _2283_/X sky130_fd_sc_hd__o31a_1
XFILLER_69_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1998_ _1998_/A vssd1 vssd1 vccd1 vccd1 _1999_/A sky130_fd_sc_hd__inv_2
X_2619_ _2848_/A _2912_/B _2619_/C _2619_/D vssd1 vssd1 vccd1 vccd1 _2619_/X sky130_fd_sc_hd__or4_2
XFILLER_18_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2970_ _1696_/A _3268_/Q _2959_/X _2969_/X vssd1 vssd1 vccd1 vccd1 _3267_/D sky130_fd_sc_hd__o211a_1
X_1921_ _1916_/X _1920_/Y _1907_/X vssd1 vssd1 vccd1 vccd1 _3001_/D sky130_fd_sc_hd__a21oi_1
X_1852_ _2995_/Q _2773_/A _1783_/X _2994_/Q vssd1 vssd1 vccd1 vccd1 _1852_/Y sky130_fd_sc_hd__a22oi_1
X_1783_ _2055_/A vssd1 vssd1 vccd1 vccd1 _1783_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3453_ _3453_/A _1624_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
X_2404_ _3095_/Q _2403_/X _2386_/X _3094_/Q vssd1 vssd1 vccd1 vccd1 _2404_/Y sky130_fd_sc_hd__a22oi_1
X_3384_ _3384_/A _1585_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2335_ _2362_/A vssd1 vssd1 vccd1 vccd1 _2335_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2266_ _2575_/B _2264_/Y _2265_/X vssd1 vssd1 vccd1 vccd1 _3049_/D sky130_fd_sc_hd__a21oi_1
X_2197_ _2194_/Y _2196_/Y _2185_/X vssd1 vssd1 vccd1 vccd1 _3036_/D sky130_fd_sc_hd__a21oi_1
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3466__92 vssd1 vssd1 vccd1 vccd1 _3466__92/HI _3466_/A sky130_fd_sc_hd__conb_1
XFILLER_31_306 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_75 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3394__36 vssd1 vssd1 vccd1 vccd1 _3394__36/HI _3394_/A sky130_fd_sc_hd__conb_1
XANTENNA_7 _2457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2120_ _3023_/Q _2097_/X _2102_/X _3022_/Q vssd1 vssd1 vccd1 vccd1 _2120_/Y sky130_fd_sc_hd__a22oi_1
Xclkbuf_leaf_23_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3242_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2051_ _3012_/Q _2050_/X _1994_/X _3011_/Q vssd1 vssd1 vccd1 vccd1 _2051_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2953_ _1714_/X _3261_/Q _2946_/X _2952_/X vssd1 vssd1 vccd1 vccd1 _3260_/D sky130_fd_sc_hd__o211a_1
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1904_ _2500_/B _2728_/B vssd1 vssd1 vccd1 vccd1 _1904_/Y sky130_fd_sc_hd__nand2_1
X_2884_ _2286_/X _2883_/Y _1679_/A vssd1 vssd1 vccd1 vccd1 _3231_/D sky130_fd_sc_hd__a21oi_1
XFILLER_30_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1835_ _2537_/B _1850_/B _1835_/C vssd1 vssd1 vccd1 vccd1 _1838_/A sky130_fd_sc_hd__or3_1
X_1766_ _3252_/Q vssd1 vssd1 vccd1 vccd1 _1890_/D sky130_fd_sc_hd__clkbuf_1
X_1697_ _3249_/Q vssd1 vssd1 vccd1 vccd1 _2550_/A sky130_fd_sc_hd__inv_2
X_3436_ _3436_/A _1609_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3367_/A _1564_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2318_ _2239_/X _2317_/Y _2309_/X vssd1 vssd1 vccd1 vccd1 _3064_/D sky130_fd_sc_hd__a21oi_1
XFILLER_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2249_ _1850_/B _2894_/A _2248_/X _1812_/X vssd1 vssd1 vccd1 vccd1 _2249_/X sky130_fd_sc_hd__a31o_1
XFILLER_82_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1620_ _1624_/A vssd1 vssd1 vccd1 vccd1 _1620_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1551_ _1575_/A vssd1 vssd1 vccd1 vccd1 _1556_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3221_ _3232_/CLK _3221_/D vssd1 vssd1 vccd1 vccd1 _3221_/Q sky130_fd_sc_hd__dfxtp_1
X_3152_ _3152_/CLK _3152_/D vssd1 vssd1 vccd1 vccd1 _3152_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2103_ _3020_/Q _2097_/X _2102_/X _3019_/Q vssd1 vssd1 vccd1 vccd1 _2103_/Y sky130_fd_sc_hd__a22oi_1
X_3083_ _3086_/CLK _3083_/D vssd1 vssd1 vccd1 vccd1 _3083_/Q sky130_fd_sc_hd__dfxtp_1
X_2034_ _2085_/B _2061_/C _2035_/B _2034_/D vssd1 vssd1 vccd1 vccd1 _2036_/A sky130_fd_sc_hd__and4b_1
XFILLER_22_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2936_ _2936_/A vssd1 vssd1 vccd1 vccd1 _3253_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2867_ _2867_/A vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__clkbuf_2
X_1818_ _1818_/A _1818_/B vssd1 vssd1 vccd1 vccd1 _2477_/B sky130_fd_sc_hd__nand2_1
X_2798_ _2796_/Y _2797_/Y _2794_/X vssd1 vssd1 vccd1 vccd1 _3201_/D sky130_fd_sc_hd__a21oi_1
X_1749_ _2901_/A _1739_/Y _2623_/C _1748_/X vssd1 vssd1 vccd1 vccd1 _1749_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_77_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3419_ _3419_/A _1542_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3436__62 vssd1 vssd1 vccd1 vccd1 _3436__62/HI _3436_/A sky130_fd_sc_hd__conb_1
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_95 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2721_ _2471_/X _2720_/Y _2665_/X vssd1 vssd1 vccd1 vccd1 _3181_/D sky130_fd_sc_hd__a21oi_1
X_2652_ _2801_/B _2651_/Y _2649_/X vssd1 vssd1 vccd1 vccd1 _3162_/D sky130_fd_sc_hd__a21oi_1
XFILLER_66_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1603_ _1605_/A vssd1 vssd1 vccd1 vccd1 _1603_/Y sky130_fd_sc_hd__inv_2
X_2583_ _2583_/A _2583_/B vssd1 vssd1 vccd1 vccd1 _2584_/B sky130_fd_sc_hd__nor2_1
X_3204_ _3230_/CLK _3204_/D vssd1 vssd1 vccd1 vccd1 _3204_/Q sky130_fd_sc_hd__dfxtp_1
X_3135_ _3168_/CLK _3135_/D vssd1 vssd1 vccd1 vccd1 _3135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3066_ _3070_/CLK _3066_/D vssd1 vssd1 vccd1 vccd1 _3066_/Q sky130_fd_sc_hd__dfxtp_1
X_2017_ _2826_/A vssd1 vssd1 vccd1 vccd1 _2017_/X sky130_fd_sc_hd__buf_2
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2919_ _2941_/S _3243_/Q vssd1 vssd1 vccd1 vccd1 _2919_/X sky130_fd_sc_hd__or2_1
XFILLER_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_504 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2704_ _3177_/Q _2704_/B vssd1 vssd1 vccd1 vccd1 _2704_/Y sky130_fd_sc_hd__nor2_1
X_2635_ _2829_/A vssd1 vssd1 vccd1 vccd1 _2635_/X sky130_fd_sc_hd__clkbuf_2
X_2566_ _2710_/B _2566_/B _2566_/C vssd1 vssd1 vccd1 vccd1 _2716_/B sky130_fd_sc_hd__nand3_2
X_2497_ _2497_/A vssd1 vssd1 vccd1 vccd1 _2638_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3118_ _3253_/CLK _3118_/D vssd1 vssd1 vccd1 vccd1 _3417_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3049_ _3062_/CLK _3049_/D vssd1 vssd1 vccd1 vccd1 _3049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2420_ _1993_/Y _2419_/Y _2416_/X vssd1 vssd1 vccd1 vccd1 _3101_/D sky130_fd_sc_hd__a21oi_1
X_2351_ _2351_/A vssd1 vssd1 vccd1 vccd1 _2351_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2282_ _2280_/X _2281_/Y _2265_/X vssd1 vssd1 vccd1 vccd1 _3052_/D sky130_fd_sc_hd__a21oi_1
XFILLER_69_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_326 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1997_ _2681_/A _1997_/B vssd1 vssd1 vccd1 vccd1 _1997_/Y sky130_fd_sc_hd__nor2_1
X_2618_ _1956_/X _2617_/Y _2600_/X vssd1 vssd1 vccd1 vccd1 _3152_/D sky130_fd_sc_hd__a21oi_1
X_2549_ _2546_/X _2547_/X _2548_/X vssd1 vssd1 vccd1 vccd1 _3131_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_470 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1920_ _3001_/Q _1919_/X _1874_/X _3000_/Q vssd1 vssd1 vccd1 vccd1 _1920_/Y sky130_fd_sc_hd__a22oi_1
X_1851_ _2756_/A _1851_/B _2905_/D vssd1 vssd1 vccd1 vccd1 _2801_/B sky130_fd_sc_hd__or3_4
X_1782_ _2101_/A vssd1 vssd1 vccd1 vccd1 _2055_/A sky130_fd_sc_hd__clkbuf_2
X_3452_ _3452_/A _1622_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
X_3383_ _3383_/A _1584_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
X_2403_ _2432_/A vssd1 vssd1 vccd1 vccd1 _2403_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2334_ _3071_/Q _2324_/X _2327_/X _3070_/Q vssd1 vssd1 vccd1 vccd1 _2334_/Y sky130_fd_sc_hd__a22oi_1
X_2265_ _2294_/A vssd1 vssd1 vccd1 vccd1 _2265_/X sky130_fd_sc_hd__clkbuf_2
X_2196_ _3036_/Q _2189_/X _2195_/X _3035_/Q vssd1 vssd1 vccd1 vccd1 _2196_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_37_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_8 _2941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2050_ _2132_/A vssd1 vssd1 vccd1 vccd1 _2050_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2952_ _2960_/A _3260_/Q vssd1 vssd1 vccd1 vccd1 _2952_/X sky130_fd_sc_hd__or2_1
X_1903_ _1903_/A vssd1 vssd1 vccd1 vccd1 _2728_/B sky130_fd_sc_hd__buf_2
X_2883_ _3231_/Q _2019_/X _2874_/X _3230_/Q vssd1 vssd1 vccd1 vccd1 _2883_/Y sky130_fd_sc_hd__a22oi_1
X_1834_ _1834_/A _1959_/A vssd1 vssd1 vccd1 vccd1 _1850_/B sky130_fd_sc_hd__or2b_1
X_1765_ _2003_/A vssd1 vssd1 vccd1 vccd1 _1765_/X sky130_fd_sc_hd__clkbuf_2
X_3435_ _3435_/A _1608_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
X_1696_ _1696_/A vssd1 vssd1 vccd1 vccd1 _1696_/X sky130_fd_sc_hd__clkbuf_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _3366_/A _1562_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _3064_/Q _2311_/X _2314_/X _3063_/Q vssd1 vssd1 vccd1 vccd1 _2317_/Y sky130_fd_sc_hd__a22oi_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _2248_/A _2248_/B _2248_/C vssd1 vssd1 vccd1 vccd1 _2248_/X sky130_fd_sc_hd__and3_2
X_2179_ _1818_/A _2583_/B _2007_/Y vssd1 vssd1 vccd1 vccd1 _2180_/B sky130_fd_sc_hd__a21o_1
XFILLER_65_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1550_ input1/X vssd1 vssd1 vccd1 vccd1 _1575_/A sky130_fd_sc_hd__clkbuf_2
X_3220_ _3234_/CLK _3220_/D vssd1 vssd1 vccd1 vccd1 _3220_/Q sky130_fd_sc_hd__dfxtp_1
X_3151_ _3154_/CLK _3151_/D vssd1 vssd1 vccd1 vccd1 _3151_/Q sky130_fd_sc_hd__dfxtp_1
X_2102_ _2227_/A vssd1 vssd1 vccd1 vccd1 _2102_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3082_ _3082_/CLK _3082_/D vssd1 vssd1 vccd1 vccd1 _3082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2033_ _2686_/A vssd1 vssd1 vccd1 vccd1 _2280_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2935_ _3406_/A _2935_/B vssd1 vssd1 vccd1 vccd1 _2936_/A sky130_fd_sc_hd__and2_1
X_2866_ _3224_/Q _2853_/X _2859_/X _3223_/Q vssd1 vssd1 vccd1 vccd1 _2866_/Y sky130_fd_sc_hd__a22oi_1
X_1817_ _2094_/B _1817_/B vssd1 vssd1 vccd1 vccd1 _1818_/B sky130_fd_sc_hd__nand2_1
X_2797_ _3201_/Q _2725_/X _2783_/X _3200_/Q vssd1 vssd1 vccd1 vccd1 _2797_/Y sky130_fd_sc_hd__a22oi_1
X_1748_ _2500_/A vssd1 vssd1 vccd1 vccd1 _1748_/X sky130_fd_sc_hd__buf_4
X_1679_ _1679_/A _1679_/B _1684_/C vssd1 vssd1 vccd1 vccd1 _2982_/D sky130_fd_sc_hd__nor3_1
X_3418_ _3418_/A _1541_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3451__77 vssd1 vssd1 vccd1 vccd1 _3451__77/HI _3451_/A sky130_fd_sc_hd__conb_1
XFILLER_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_262 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2720_ _3181_/Q _2653_/X _2656_/X _3180_/Q vssd1 vssd1 vccd1 vccd1 _2720_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2651_ _3162_/Q _2635_/X _2642_/X _3161_/Q vssd1 vssd1 vccd1 vccd1 _2651_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_8_163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1602_ _1605_/A vssd1 vssd1 vccd1 vccd1 _1602_/Y sky130_fd_sc_hd__inv_2
X_2582_ _2041_/X _2581_/Y _2572_/X vssd1 vssd1 vccd1 vccd1 _3140_/D sky130_fd_sc_hd__a21oi_1
XFILLER_59_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3203_ _3233_/CLK _3203_/D vssd1 vssd1 vccd1 vccd1 _3203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3134_ _3152_/CLK _3134_/D vssd1 vssd1 vccd1 vccd1 _3134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3065_ _3070_/CLK _3065_/D vssd1 vssd1 vccd1 vccd1 _3065_/Q sky130_fd_sc_hd__dfxtp_1
X_2016_ _2728_/A vssd1 vssd1 vccd1 vccd1 _2826_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2918_ _2918_/A vssd1 vssd1 vccd1 vccd1 _3242_/D sky130_fd_sc_hd__clkbuf_1
X_2849_ _3217_/Q _2829_/X _2832_/X _3216_/Q vssd1 vssd1 vccd1 vccd1 _2849_/Y sky130_fd_sc_hd__a22oi_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_398 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2703_ _2500_/D _2701_/X _2596_/Y _2702_/Y _2280_/A vssd1 vssd1 vccd1 vccd1 _2703_/X
+ sky130_fd_sc_hd__a32o_1
X_2634_ _2634_/A vssd1 vssd1 vccd1 vccd1 _2829_/A sky130_fd_sc_hd__clkbuf_2
X_2565_ _3135_/Q _2512_/X _2564_/X _2517_/X vssd1 vssd1 vccd1 vccd1 _3135_/D sky130_fd_sc_hd__o211a_1
X_2496_ _2496_/A vssd1 vssd1 vccd1 vccd1 _3122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3117_ _3253_/CLK _3117_/D vssd1 vssd1 vccd1 vccd1 _3117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3048_ _3062_/CLK _3048_/D vssd1 vssd1 vccd1 vccd1 _3048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3421__47 vssd1 vssd1 vccd1 vccd1 _3421__47/HI _3421_/A sky130_fd_sc_hd__conb_1
XFILLER_23_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3062_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2350_ _2171_/Y _2348_/Y _2349_/X vssd1 vssd1 vccd1 vccd1 _3076_/D sky130_fd_sc_hd__a21oi_1
X_2281_ _3052_/Q _2271_/X _2277_/X _3051_/Q vssd1 vssd1 vccd1 vccd1 _2281_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_346 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1996_ _1993_/Y _1995_/Y _1976_/X vssd1 vssd1 vccd1 vccd1 _3007_/D sky130_fd_sc_hd__a21oi_1
XFILLER_20_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2617_ _3152_/Q _2606_/X _2611_/X _3151_/Q vssd1 vssd1 vccd1 vccd1 _2617_/Y sky130_fd_sc_hd__a22oi_1
X_2548_ _3131_/Q _2507_/X _2483_/X _3130_/Q _2939_/B vssd1 vssd1 vccd1 vccd1 _2548_/X
+ sky130_fd_sc_hd__o221a_1
X_2479_ _2621_/A vssd1 vssd1 vccd1 vccd1 _2479_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_408 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_110 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1850_ _2538_/A _1850_/B vssd1 vssd1 vccd1 vccd1 _2905_/D sky130_fd_sc_hd__nand2_2
X_1781_ _2250_/A vssd1 vssd1 vccd1 vccd1 _2101_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3451_ _3451_/A _1620_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3382_ _3382_/A _1583_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
X_2402_ _2064_/X _2400_/Y _2401_/X vssd1 vssd1 vccd1 vccd1 _3094_/D sky130_fd_sc_hd__a21oi_1
X_2333_ _2207_/Y _2332_/Y _2322_/X vssd1 vssd1 vccd1 vccd1 _3070_/D sky130_fd_sc_hd__a21oi_1
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2264_ _3049_/Q _2244_/X _2252_/X _3048_/Q vssd1 vssd1 vccd1 vccd1 _2264_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2195_ _2227_/A vssd1 vssd1 vccd1 vccd1 _2195_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_400 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1979_ _2026_/B _1979_/B vssd1 vssd1 vccd1 vccd1 _2912_/C sky130_fd_sc_hd__nor2_4
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 _3248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3457__83 vssd1 vssd1 vccd1 vccd1 _3457__83/HI _3457_/A sky130_fd_sc_hd__conb_1
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2951_ _1714_/X _3260_/Q _2946_/X _2950_/X vssd1 vssd1 vccd1 vccd1 _3259_/D sky130_fd_sc_hd__o211a_1
XFILLER_62_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_32_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3185_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1902_ _1913_/B _1913_/C _1893_/B vssd1 vssd1 vccd1 vccd1 _1903_/A sky130_fd_sc_hd__or3b_1
X_2882_ _2286_/X _2881_/Y _1679_/A vssd1 vssd1 vccd1 vccd1 _3230_/D sky130_fd_sc_hd__a21oi_1
XFILLER_30_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1833_ _2085_/B vssd1 vssd1 vccd1 vccd1 _2537_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3385__27 vssd1 vssd1 vccd1 vccd1 _3385__27/HI _3385_/A sky130_fd_sc_hd__conb_1
X_1764_ _2034_/D _2061_/D vssd1 vssd1 vccd1 vccd1 _2003_/A sky130_fd_sc_hd__nor2_2
X_3434_ _3434_/A _1607_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
X_1695_ _2584_/A vssd1 vssd1 vccd1 vccd1 _1696_/A sky130_fd_sc_hd__buf_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _3365_/A _1561_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _2243_/Y _2315_/Y _2309_/X vssd1 vssd1 vccd1 vccd1 _3063_/D sky130_fd_sc_hd__a21oi_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _2128_/A _2004_/A _2566_/C vssd1 vssd1 vccd1 vccd1 _2248_/C sky130_fd_sc_hd__o21a_1
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2178_ _2178_/A vssd1 vssd1 vccd1 vccd1 _2583_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_53_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3150_ _3253_/CLK _3150_/D vssd1 vssd1 vccd1 vccd1 _3150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2101_ _2101_/A vssd1 vssd1 vccd1 vccd1 _2227_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3081_ _3082_/CLK _3081_/D vssd1 vssd1 vccd1 vccd1 _3081_/Q sky130_fd_sc_hd__dfxtp_1
X_2032_ _2032_/A vssd1 vssd1 vccd1 vccd1 _2686_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_411 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2934_ _2934_/A vssd1 vssd1 vccd1 vccd1 _3252_/D sky130_fd_sc_hd__clkbuf_1
X_2865_ _2810_/Y _2864_/Y _2846_/X vssd1 vssd1 vccd1 vccd1 _3223_/D sky130_fd_sc_hd__a21oi_1
X_1816_ _1936_/A _1924_/B vssd1 vssd1 vccd1 vccd1 _2094_/B sky130_fd_sc_hd__nor2b_2
XFILLER_7_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2796_ _2532_/A _2570_/C _2164_/X _2275_/X vssd1 vssd1 vccd1 vccd1 _2796_/Y sky130_fd_sc_hd__o31ai_4
X_1747_ _1897_/A vssd1 vssd1 vccd1 vccd1 _2500_/A sky130_fd_sc_hd__clkbuf_2
X_1678_ _3410_/A _3411_/A _3412_/A vssd1 vssd1 vccd1 vccd1 _1684_/C sky130_fd_sc_hd__and3_1
X_3417_ _3417_/A _1540_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_75 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3427__53 vssd1 vssd1 vccd1 vccd1 _3427__53/HI _3427_/A sky130_fd_sc_hd__conb_1
XFILLER_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2650_ _2619_/X _2647_/Y _2649_/X vssd1 vssd1 vccd1 vccd1 _3161_/D sky130_fd_sc_hd__a21oi_1
X_1601_ _1605_/A vssd1 vssd1 vccd1 vccd1 _1601_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2581_ _3140_/Q _2580_/X _2559_/X _3139_/Q vssd1 vssd1 vccd1 vccd1 _2581_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_4_381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3202_ _3233_/CLK _3202_/D vssd1 vssd1 vccd1 vccd1 _3202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3133_ _3152_/CLK _3133_/D vssd1 vssd1 vccd1 vccd1 _3133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3064_ _3070_/CLK _3064_/D vssd1 vssd1 vccd1 vccd1 _3064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2015_ _2015_/A _2567_/C _2825_/B vssd1 vssd1 vccd1 vccd1 _2015_/X sky130_fd_sc_hd__or3_1
XFILLER_23_414 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2917_ _2959_/A _2917_/B _2917_/C vssd1 vssd1 vccd1 vccd1 _2918_/A sky130_fd_sc_hd__and3_1
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2848_ _2848_/A _2848_/B _2915_/A _2848_/D vssd1 vssd1 vccd1 vccd1 _2848_/X sky130_fd_sc_hd__or4_1
X_2779_ _2007_/Y _2268_/A _2474_/B _1835_/C _2538_/A vssd1 vssd1 vccd1 vccd1 _2779_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_344 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2702_ _3176_/Q vssd1 vssd1 vccd1 vccd1 _2702_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2633_ _2498_/X _2630_/X _2631_/X _2632_/X vssd1 vssd1 vccd1 vccd1 _3156_/D sky130_fd_sc_hd__o211a_1
X_2564_ _2562_/Y _2563_/X _2638_/A vssd1 vssd1 vccd1 vccd1 _2564_/X sky130_fd_sc_hd__a21o_1
X_2495_ _2524_/A _2495_/B _2495_/C vssd1 vssd1 vccd1 vccd1 _2496_/A sky130_fd_sc_hd__and3_1
X_3116_ _3116_/CLK _3116_/D vssd1 vssd1 vccd1 vccd1 _3116_/Q sky130_fd_sc_hd__dfxtp_1
X_3047_ _3062_/CLK _3047_/D vssd1 vssd1 vccd1 vccd1 _3047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2280_ _2280_/A _2280_/B vssd1 vssd1 vccd1 vccd1 _2280_/X sky130_fd_sc_hd__or2_1
XFILLER_77_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1995_ _3007_/Q _1986_/X _1994_/X _3006_/Q vssd1 vssd1 vccd1 vccd1 _1995_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2616_ _2498_/X _2614_/X _2615_/X _2517_/X vssd1 vssd1 vccd1 vccd1 _3151_/D sky130_fd_sc_hd__o211a_1
X_2547_ _2547_/A _2788_/B _2547_/C _2667_/D vssd1 vssd1 vccd1 vccd1 _2547_/X sky130_fd_sc_hd__or4_1
X_2478_ _3120_/Q _2460_/X _2463_/X _3119_/Q vssd1 vssd1 vccd1 vccd1 _2478_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_18_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1780_ _2481_/A _3404_/A vssd1 vssd1 vccd1 vccd1 _2250_/A sky130_fd_sc_hd__and2_1
X_3450_ _3450_/A _1617_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
X_3381_ _3381_/A _1580_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
X_2401_ _2443_/A vssd1 vssd1 vccd1 vccd1 _2401_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2332_ _3070_/Q _2324_/X _2327_/X _3069_/Q vssd1 vssd1 vccd1 vccd1 _2332_/Y sky130_fd_sc_hd__a22oi_1
X_2263_ _2567_/C _2716_/A _2693_/D vssd1 vssd1 vccd1 vccd1 _2575_/B sky130_fd_sc_hd__or3_4
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2194_ _1991_/B _1991_/D _2193_/X _2165_/X vssd1 vssd1 vccd1 vccd1 _2194_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_65_431 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1978_ _2756_/A vssd1 vssd1 vccd1 vccd1 _2912_/B sky130_fd_sc_hd__buf_2
XFILLER_0_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3105_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2950_ _2960_/A _3259_/Q vssd1 vssd1 vccd1 vccd1 _2950_/X sky130_fd_sc_hd__or2_1
XFILLER_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1901_ _1899_/Y _1900_/Y _1853_/X vssd1 vssd1 vccd1 vccd1 _2999_/D sky130_fd_sc_hd__a21oi_1
X_2881_ _3230_/Q _2871_/X _2874_/X _3229_/Q vssd1 vssd1 vccd1 vccd1 _2881_/Y sky130_fd_sc_hd__a22oi_1
X_1832_ _1998_/A vssd1 vssd1 vccd1 vccd1 _2085_/B sky130_fd_sc_hd__clkbuf_1
X_1763_ _2058_/A vssd1 vssd1 vccd1 vccd1 _2061_/D sky130_fd_sc_hd__clkbuf_2
X_1694_ _2032_/A vssd1 vssd1 vccd1 vccd1 _2584_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3433_ _3433_/A _1654_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3364_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _3063_/Q _2311_/X _2314_/X _3062_/Q vssd1 vssd1 vccd1 vccd1 _2315_/Y sky130_fd_sc_hd__a22oi_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _2243_/Y _2245_/Y _2241_/X vssd1 vssd1 vccd1 vccd1 _3045_/D sky130_fd_sc_hd__a21oi_1
XFILLER_65_250 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2177_ _2175_/X _2176_/Y _2155_/X vssd1 vssd1 vccd1 vccd1 _3033_/D sky130_fd_sc_hd__a21oi_1
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2100_ _2780_/A _1819_/X _2905_/B _2492_/B _1748_/X vssd1 vssd1 vccd1 vccd1 _2100_/Y
+ sky130_fd_sc_hd__o41ai_4
X_3080_ _3080_/CLK _3080_/D vssd1 vssd1 vccd1 vccd1 _3080_/Q sky130_fd_sc_hd__dfxtp_1
X_2031_ _2029_/Y _2030_/Y _1976_/X vssd1 vssd1 vccd1 vccd1 _3010_/D sky130_fd_sc_hd__a21oi_1
XFILLER_35_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2933_ _3405_/A _2935_/B vssd1 vssd1 vccd1 vccd1 _2934_/A sky130_fd_sc_hd__and2_1
XFILLER_50_437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2864_ _3223_/Q _2853_/X _2859_/X _3222_/Q vssd1 vssd1 vccd1 vccd1 _2864_/Y sky130_fd_sc_hd__a22oi_1
X_1815_ _1813_/X _1814_/Y _1672_/B vssd1 vssd1 vccd1 vccd1 _2993_/D sky130_fd_sc_hd__a21oi_1
X_2795_ _2792_/Y _2793_/Y _2794_/X vssd1 vssd1 vccd1 vccd1 _3200_/D sky130_fd_sc_hd__a21oi_1
X_1746_ _2538_/A vssd1 vssd1 vccd1 vccd1 _1897_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1677_ _3410_/A _3411_/A _3412_/A vssd1 vssd1 vccd1 vccd1 _1679_/B sky130_fd_sc_hd__a21oi_1
X_3416_ _3416_/A _1539_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ _2226_/Y _2228_/Y _2214_/X vssd1 vssd1 vccd1 vccd1 _3041_/D sky130_fd_sc_hd__a21oi_1
XFILLER_26_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3442__68 vssd1 vssd1 vccd1 vccd1 _3442__68/HI _3442_/A sky130_fd_sc_hd__conb_1
XFILLER_40_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1600_ _1606_/A vssd1 vssd1 vccd1 vccd1 _1605_/A sky130_fd_sc_hd__clkbuf_4
X_2580_ _2606_/A vssd1 vssd1 vccd1 vccd1 _2580_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3201_ _3233_/CLK _3201_/D vssd1 vssd1 vccd1 vccd1 _3201_/Q sky130_fd_sc_hd__dfxtp_1
X_3132_ _3157_/CLK _3132_/D vssd1 vssd1 vccd1 vccd1 _3132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3063_ _3070_/CLK _3063_/D vssd1 vssd1 vccd1 vccd1 _3063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2014_ _2067_/A _2268_/B _2129_/B _2748_/A vssd1 vssd1 vccd1 vccd1 _2825_/B sky130_fd_sc_hd__a22o_1
XFILLER_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2916_ _3242_/Q _2687_/X _2483_/A _3241_/Q vssd1 vssd1 vccd1 vccd1 _2917_/C sky130_fd_sc_hd__o22a_1
XFILLER_50_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2847_ _2217_/Y _2845_/Y _2846_/X vssd1 vssd1 vccd1 vccd1 _3216_/D sky130_fd_sc_hd__a21oi_1
X_2778_ _2788_/A _2778_/B vssd1 vssd1 vccd1 vccd1 _2778_/X sky130_fd_sc_hd__or2_1
X_1729_ _3251_/Q vssd1 vssd1 vccd1 vccd1 _1888_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2701_ _2500_/B _1765_/X _2045_/C _2583_/B _2500_/C vssd1 vssd1 vccd1 vccd1 _2701_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2632_ _2843_/A vssd1 vssd1 vccd1 vccd1 _2632_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2563_ _2826_/A _3134_/Q vssd1 vssd1 vccd1 vccd1 _2563_/X sky130_fd_sc_hd__or2_1
X_2494_ _3122_/Q _2511_/A _2493_/X _3121_/Q vssd1 vssd1 vccd1 vccd1 _2495_/C sky130_fd_sc_hd__o22a_1
XFILLER_4_72 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3115_ _3116_/CLK _3115_/D vssd1 vssd1 vccd1 vccd1 _3115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3046_ _3062_/CLK _3046_/D vssd1 vssd1 vccd1 vccd1 _3046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_440 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3248_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1994_ _2055_/A vssd1 vssd1 vccd1 vccd1 _1994_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2615_ _3151_/Q _2660_/B vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__or2_1
X_2546_ _2905_/B _2905_/C _2546_/C vssd1 vssd1 vccd1 vccd1 _2546_/X sky130_fd_sc_hd__or3_1
X_2477_ _2477_/A _2477_/B _2477_/C _2477_/D vssd1 vssd1 vccd1 vccd1 _2477_/X sky130_fd_sc_hd__or4_1
X_3029_ _3082_/CLK _3029_/D vssd1 vssd1 vccd1 vccd1 _3029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2400_ _3094_/Q _2383_/X _2386_/X _3093_/Q vssd1 vssd1 vccd1 vccd1 _2400_/Y sky130_fd_sc_hd__a22oi_1
X_3380_ _3380_/A _1579_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
X_2331_ _2212_/Y _2330_/Y _2322_/X vssd1 vssd1 vccd1 vccd1 _3069_/D sky130_fd_sc_hd__a21oi_1
XFILLER_69_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2262_ _2728_/A _2262_/B vssd1 vssd1 vccd1 vccd1 _2693_/D sky130_fd_sc_hd__nand2_2
XFILLER_69_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2193_ _2198_/A _2681_/A _2681_/B _2912_/D vssd1 vssd1 vccd1 vccd1 _2193_/X sky130_fd_sc_hd__or4_1
XFILLER_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1977_ _1972_/Y _1973_/Y _1976_/X vssd1 vssd1 vccd1 vccd1 _3005_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2529_ _3127_/Q _2527_/X _2528_/X _3126_/Q _2959_/A vssd1 vssd1 vccd1 vccd1 _2529_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1900_ _2999_/Q _1863_/X _1874_/X _2998_/Q vssd1 vssd1 vccd1 vccd1 _1900_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2880_ _2562_/Y _2879_/Y _1679_/A vssd1 vssd1 vccd1 vccd1 _3229_/D sky130_fd_sc_hd__a21oi_1
X_1831_ _2204_/A _2885_/A _2015_/A _1831_/D vssd1 vssd1 vccd1 vccd1 _1831_/X sky130_fd_sc_hd__or4_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1762_ _1924_/A vssd1 vssd1 vccd1 vccd1 _2034_/D sky130_fd_sc_hd__clkbuf_2
X_1693_ _2481_/A vssd1 vssd1 vccd1 vccd1 _2032_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3432_ _3432_/A _1605_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
X_3363_ _3363_/A _1559_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _2327_/A vssd1 vssd1 vccd1 vccd1 _2314_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _3045_/Q _2244_/X _2227_/X _3044_/Q vssd1 vssd1 vccd1 vccd1 _2245_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2176_ _3033_/Q _2159_/X _2167_/X _3032_/Q vssd1 vssd1 vccd1 vccd1 _2176_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_38_454 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3448__74 vssd1 vssd1 vccd1 vccd1 _3448__74/HI _3448_/A sky130_fd_sc_hd__conb_1
XFILLER_80_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3376__18 vssd1 vssd1 vccd1 vccd1 _3376__18/HI _3376_/A sky130_fd_sc_hd__conb_1
XFILLER_0_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_118 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3390__32 vssd1 vssd1 vccd1 vccd1 _3390__32/HI _3390_/A sky130_fd_sc_hd__conb_1
XFILLER_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2030_ _3010_/Q _1986_/X _1994_/X _3009_/Q vssd1 vssd1 vccd1 vccd1 _2030_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2932_ _2932_/A vssd1 vssd1 vccd1 vccd1 _3251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2863_ _2905_/D _2519_/C _2862_/X vssd1 vssd1 vccd1 vccd1 _3222_/D sky130_fd_sc_hd__o21a_1
X_1814_ _2993_/Q _2773_/A _1783_/X _2992_/Q vssd1 vssd1 vccd1 vccd1 _1814_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2794_ _2846_/A vssd1 vssd1 vccd1 vccd1 _2794_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1745_ _2686_/B vssd1 vssd1 vccd1 vccd1 _2623_/C sky130_fd_sc_hd__clkbuf_2
X_1676_ _2867_/A vssd1 vssd1 vccd1 vccd1 _1679_/A sky130_fd_sc_hd__clkbuf_2
X_3415_ _3415_/A _1669_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ _3041_/Q _2218_/X _2227_/X _3040_/Q vssd1 vssd1 vccd1 vccd1 _2228_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_26_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2159_ _2271_/A vssd1 vssd1 vccd1 vccd1 _2159_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_162 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3200_ _3233_/CLK _3200_/D vssd1 vssd1 vccd1 vccd1 _3200_/Q sky130_fd_sc_hd__dfxtp_1
X_3131_ _3154_/CLK _3131_/D vssd1 vssd1 vccd1 vccd1 _3131_/Q sky130_fd_sc_hd__dfxtp_1
X_3062_ _3062_/CLK _3062_/D vssd1 vssd1 vccd1 vccd1 _3062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2013_ _2013_/A _1887_/B vssd1 vssd1 vccd1 vccd1 _2567_/C sky130_fd_sc_hd__or2b_2
XFILLER_31_471 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2915_ _2915_/A _2915_/B _2915_/C _2566_/C vssd1 vssd1 vccd1 vccd1 _2917_/B sky130_fd_sc_hd__or4b_1
X_2846_ _2846_/A vssd1 vssd1 vccd1 vccd1 _2846_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2777_ _2773_/X _2775_/X _2776_/X _2708_/X vssd1 vssd1 vccd1 vccd1 _3195_/D sky130_fd_sc_hd__o211a_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1728_ _1946_/A _1947_/C _1804_/A vssd1 vssd1 vccd1 vccd1 _1968_/A sky130_fd_sc_hd__and3b_1
X_1659_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1659_/Y sky130_fd_sc_hd__inv_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2700_ _2638_/X _2698_/X _2699_/X _2632_/X vssd1 vssd1 vccd1 vccd1 _3176_/D sky130_fd_sc_hd__o211a_1
XFILLER_43_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2631_ _3156_/Q _2660_/B vssd1 vssd1 vccd1 vccd1 _2631_/X sky130_fd_sc_hd__or2_1
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2562_ _2223_/Y _1962_/X _2699_/A vssd1 vssd1 vccd1 vccd1 _2562_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2493_ _2624_/A vssd1 vssd1 vccd1 vccd1 _2493_/X sky130_fd_sc_hd__clkbuf_2
X_3114_ _3116_/CLK _3114_/D vssd1 vssd1 vccd1 vccd1 _3114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3045_ _3062_/CLK _3045_/D vssd1 vssd1 vccd1 vccd1 _3045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2829_ _2829_/A vssd1 vssd1 vccd1 vccd1 _2829_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_110 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_308 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_452 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1993_ _1997_/B _2552_/B _2471_/D _1992_/X vssd1 vssd1 vccd1 vccd1 _1993_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_60_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2614_ _1811_/Y _2513_/X _2699_/A _3150_/Q vssd1 vssd1 vccd1 vccd1 _2614_/X sky130_fd_sc_hd__o2bb2a_1
X_2545_ _2892_/B _2544_/Y _2479_/X vssd1 vssd1 vccd1 vccd1 _3130_/D sky130_fd_sc_hd__a21oi_1
X_2476_ _2547_/A _2547_/C _2667_/D vssd1 vssd1 vccd1 vccd1 _2477_/D sky130_fd_sc_hd__or3_2
XFILLER_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3028_ _3028_/CLK _3028_/D vssd1 vssd1 vccd1 vccd1 _3028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_264 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2330_ _3069_/Q _2324_/X _2327_/X _3068_/Q vssd1 vssd1 vccd1 vccd1 _2330_/Y sky130_fd_sc_hd__a22oi_1
X_2261_ _2259_/Y _2260_/Y _2241_/X vssd1 vssd1 vccd1 vccd1 _3048_/D sky130_fd_sc_hd__a21oi_1
XFILLER_2_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2192_ _2199_/B _2526_/B vssd1 vssd1 vccd1 vccd1 _2912_/D sky130_fd_sc_hd__nor2_1
XFILLER_37_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1976_ _2155_/A vssd1 vssd1 vccd1 vccd1 _1976_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2528_ _2767_/A vssd1 vssd1 vccd1 vccd1 _2528_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2459_ _1813_/X _2456_/Y _2458_/X vssd1 vssd1 vccd1 vccd1 _3115_/D sky130_fd_sc_hd__a21oi_1
XFILLER_28_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1830_ _1829_/X _1935_/A _1961_/A vssd1 vssd1 vccd1 vccd1 _1831_/D sky130_fd_sc_hd__a21o_1
X_1761_ _1834_/A vssd1 vssd1 vccd1 vccd1 _2223_/B sky130_fd_sc_hd__buf_2
X_1692_ _3403_/A vssd1 vssd1 vccd1 vccd1 _2481_/A sky130_fd_sc_hd__inv_2
X_3431_ _3431_/A _1558_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2249_/X _2312_/Y _2309_/X vssd1 vssd1 vccd1 vccd1 _3062_/D sky130_fd_sc_hd__a21oi_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _2271_/A vssd1 vssd1 vccd1 vccd1 _2244_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3028_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2175_ _2677_/A _2686_/C _2175_/C vssd1 vssd1 vccd1 vccd1 _2175_/X sky130_fd_sc_hd__or3_4
XFILLER_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3463__89 vssd1 vssd1 vccd1 vccd1 _3463__89/HI _3463_/A sky130_fd_sc_hd__conb_1
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_480 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1959_ _1959_/A _2223_/B vssd1 vssd1 vccd1 vccd1 _2046_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_422 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _2987_/Q _2935_/B vssd1 vssd1 vccd1 vccd1 _2932_/A sky130_fd_sc_hd__and2_1
X_2862_ _3222_/Q _2761_/X _2528_/X _3221_/Q _2524_/A vssd1 vssd1 vccd1 vccd1 _2862_/X
+ sky130_fd_sc_hd__o221a_1
X_1813_ _2500_/B _2075_/A _2894_/A _1811_/Y _1812_/X vssd1 vssd1 vccd1 vccd1 _1813_/X
+ sky130_fd_sc_hd__a41o_1
X_2793_ _3200_/Q _2725_/X _2783_/X _3199_/Q vssd1 vssd1 vccd1 vccd1 _2793_/Y sky130_fd_sc_hd__a22oi_1
X_1744_ _1817_/B vssd1 vssd1 vccd1 vccd1 _2686_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3414_ _3414_/A _1668_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
X_1675_ _2980_/Q _3411_/A _1674_/Y vssd1 vssd1 vccd1 vccd1 _2981_/D sky130_fd_sc_hd__o21a_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _2227_/A vssd1 vssd1 vccd1 vccd1 _2227_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2158_ _2296_/A vssd1 vssd1 vccd1 vccd1 _2271_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2089_ _2848_/D vssd1 vssd1 vccd1 vccd1 _2532_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3130_ _3154_/CLK _3130_/D vssd1 vssd1 vccd1 vccd1 _3130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_314 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3061_ _3062_/CLK _3061_/D vssd1 vssd1 vccd1 vccd1 _3061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2012_ _2012_/A vssd1 vssd1 vccd1 vccd1 _2848_/B sky130_fd_sc_hd__buf_2
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3433__59 vssd1 vssd1 vccd1 vccd1 _3433__59/HI _3433_/A sky130_fd_sc_hd__conb_1
X_2914_ _2467_/A _2667_/D _2912_/X _2913_/X vssd1 vssd1 vccd1 vccd1 _3241_/D sky130_fd_sc_hd__o31a_1
XFILLER_12_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2845_ _3216_/Q _2829_/X _2832_/X _3215_/Q vssd1 vssd1 vccd1 vccd1 _2845_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_12_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2776_ _3195_/Q _2842_/B vssd1 vssd1 vccd1 vccd1 _2776_/X sky130_fd_sc_hd__or2_1
X_1727_ _3253_/Q vssd1 vssd1 vccd1 vccd1 _1804_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1658_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1658_/Y sky130_fd_sc_hd__inv_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ _1593_/A vssd1 vssd1 vccd1 vccd1 _1589_/Y sky130_fd_sc_hd__inv_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3259_ _3270_/CLK _3259_/D vssd1 vssd1 vccd1 vccd1 _3259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2630_ _2973_/A _3155_/Q _1739_/Y _2500_/Y vssd1 vssd1 vccd1 vccd1 _2630_/X sky130_fd_sc_hd__o22a_1
X_2561_ _1956_/X _2560_/Y _2479_/X vssd1 vssd1 vccd1 vccd1 _3134_/D sky130_fd_sc_hd__a21oi_1
X_2492_ _2686_/A _2492_/B _2492_/C _2519_/D vssd1 vssd1 vccd1 vccd1 _2495_/B sky130_fd_sc_hd__or4_1
XFILLER_4_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3113_ _3113_/CLK _3113_/D vssd1 vssd1 vccd1 vccd1 _3113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3044_ _3070_/CLK _3044_/D vssd1 vssd1 vccd1 vccd1 _3044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2828_ _3210_/Q _2512_/X _2827_/X _2708_/X vssd1 vssd1 vccd1 vccd1 _3210_/D sky130_fd_sc_hd__o211a_1
X_2759_ _2170_/A _2583_/B _1880_/X _1857_/A _1897_/A vssd1 vssd1 vccd1 vccd1 _2760_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1992_ _2752_/A vssd1 vssd1 vccd1 vccd1 _1992_/X sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_35_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3157_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2613_ _1985_/Y _2612_/Y _2600_/X vssd1 vssd1 vccd1 vccd1 _3150_/D sky130_fd_sc_hd__a21oi_1
X_2544_ _3130_/Q _2460_/X _2463_/X _3129_/Q vssd1 vssd1 vccd1 vccd1 _2544_/Y sky130_fd_sc_hd__a22oi_1
X_2475_ _1739_/B _1889_/X _2481_/A vssd1 vssd1 vccd1 vccd1 _2667_/D sky130_fd_sc_hd__a21o_1
XFILLER_55_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3027_ _3028_/CLK _3027_/D vssd1 vssd1 vccd1 vccd1 _3027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3469__95 vssd1 vssd1 vccd1 vccd1 _3469__95/HI _3469_/A sky130_fd_sc_hd__conb_1
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3397__39 vssd1 vssd1 vccd1 vccd1 _3397__39/HI _3397_/A sky130_fd_sc_hd__conb_1
XFILLER_24_71 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_276 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2260_ _3048_/Q _2244_/X _2252_/X _3047_/Q vssd1 vssd1 vccd1 vccd1 _2260_/Y sky130_fd_sc_hd__a22oi_1
X_2191_ _2188_/X _2190_/Y _2185_/X vssd1 vssd1 vccd1 vccd1 _3035_/D sky130_fd_sc_hd__a21oi_1
XFILLER_1_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1975_ _2457_/A vssd1 vssd1 vccd1 vccd1 _2155_/A sky130_fd_sc_hd__clkbuf_2
X_2527_ _2761_/A vssd1 vssd1 vccd1 vccd1 _2527_/X sky130_fd_sc_hd__clkbuf_2
X_2458_ _2621_/A vssd1 vssd1 vccd1 vccd1 _2458_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2389_ _3090_/Q _2383_/X _2386_/X _3089_/Q vssd1 vssd1 vccd1 vccd1 _2389_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1760_ _1960_/D vssd1 vssd1 vccd1 vccd1 _1834_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1691_ _3416_/A _2929_/C _3247_/D vssd1 vssd1 vccd1 vccd1 _2986_/D sky130_fd_sc_hd__o21a_1
X_3430_ _3430_/A _1556_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2312_ _3062_/Q _2311_/X _2300_/X _3061_/Q vssd1 vssd1 vccd1 vccd1 _2312_/Y sky130_fd_sc_hd__a22oi_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2243_ _2519_/C _2064_/C _1898_/X vssd1 vssd1 vccd1 vccd1 _2243_/Y sky130_fd_sc_hd__o21ai_2
X_2174_ _2738_/A vssd1 vssd1 vccd1 vccd1 _2677_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1958_ _1956_/X _1957_/Y _1907_/X vssd1 vssd1 vccd1 vccd1 _3004_/D sky130_fd_sc_hd__a21oi_1
X_1889_ _2267_/B vssd1 vssd1 vccd1 vccd1 _1889_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3439__65 vssd1 vssd1 vccd1 vccd1 _3439__65/HI _3439_/A sky130_fd_sc_hd__conb_1
XFILLER_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2930_ _2930_/A vssd1 vssd1 vccd1 vccd1 _3248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2861_ _2243_/Y _2860_/Y _2846_/X vssd1 vssd1 vccd1 vccd1 _3221_/D sky130_fd_sc_hd__a21oi_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2792_ _2912_/A _2888_/A _2716_/B _2275_/X vssd1 vssd1 vccd1 vccd1 _2792_/Y sky130_fd_sc_hd__o31ai_4
X_1812_ _2765_/B vssd1 vssd1 vccd1 vccd1 _1812_/X sky130_fd_sc_hd__clkbuf_2
X_1743_ _2061_/C _1960_/D _1960_/B vssd1 vssd1 vccd1 vccd1 _1817_/B sky130_fd_sc_hd__and3b_1
XFILLER_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1674_ _3410_/A _3411_/A _1681_/A vssd1 vssd1 vccd1 vccd1 _1674_/Y sky130_fd_sc_hd__a21oi_1
X_3413_ _3413_/A _1667_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
X_3381__23 vssd1 vssd1 vccd1 vccd1 _3381__23/HI _3381_/A sky130_fd_sc_hd__conb_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _2222_/X _2224_/X _2526_/A vssd1 vssd1 vccd1 vccd1 _2226_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2157_ _2584_/A _2157_/B _2157_/C vssd1 vssd1 vccd1 vccd1 _2157_/X sky130_fd_sc_hd__or3_2
X_2088_ _2248_/A _2248_/B vssd1 vssd1 vccd1 vccd1 _2848_/D sky130_fd_sc_hd__nand2_1
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3060_ _3062_/CLK _3060_/D vssd1 vssd1 vccd1 vccd1 _3060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2011_ _2009_/X _2010_/Y _1976_/X vssd1 vssd1 vccd1 vccd1 _3008_/D sky130_fd_sc_hd__a21oi_1
XFILLER_67_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2913_ _3241_/Q _2542_/B _2493_/X _3240_/Q _2929_/B vssd1 vssd1 vccd1 vccd1 _2913_/X
+ sky130_fd_sc_hd__o221a_1
X_2844_ _2773_/X _2841_/X _2842_/X _2843_/X vssd1 vssd1 vccd1 vccd1 _3215_/D sky130_fd_sc_hd__o211a_1
X_2775_ _2912_/A _2888_/A _2774_/X _3194_/Q _1705_/A vssd1 vssd1 vccd1 vccd1 _2775_/X
+ sky130_fd_sc_hd__o32a_1
X_1726_ _1794_/A vssd1 vssd1 vccd1 vccd1 _1947_/C sky130_fd_sc_hd__clkbuf_1
X_1657_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1657_/Y sky130_fd_sc_hd__inv_2
X_1588_ _1606_/A vssd1 vssd1 vccd1 vccd1 _1593_/A sky130_fd_sc_hd__buf_6
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3258_ _3270_/CLK _3258_/D vssd1 vssd1 vccd1 vccd1 _3258_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2209_ _2207_/Y _2208_/Y _2185_/X vssd1 vssd1 vccd1 vccd1 _3038_/D sky130_fd_sc_hd__a21oi_1
XFILLER_73_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3189_ _3269_/CLK _3189_/D vssd1 vssd1 vccd1 vccd1 _3189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2560_ _3134_/Q _2556_/X _2559_/X _3133_/Q vssd1 vssd1 vccd1 vccd1 _2560_/Y sky130_fd_sc_hd__a22oi_1
X_2491_ _1963_/A _2128_/A _2067_/A _2094_/B _2788_/B vssd1 vssd1 vccd1 vccd1 _2519_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_4_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3112_ _3113_/CLK _3112_/D vssd1 vssd1 vccd1 vccd1 _3112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3043_ _3070_/CLK _3043_/D vssd1 vssd1 vccd1 vccd1 _3043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2827_ _2825_/X _2826_/X _2638_/A vssd1 vssd1 vccd1 vccd1 _2827_/X sky130_fd_sc_hd__a21o_1
X_2758_ _3191_/Q _2512_/X _2757_/X _2708_/X vssd1 vssd1 vccd1 vccd1 _3191_/D sky130_fd_sc_hd__o211a_1
X_1709_ _1696_/X _3406_/A _1700_/X _1708_/X vssd1 vssd1 vccd1 vccd1 _2988_/D sky130_fd_sc_hd__o211a_1
X_2689_ _2689_/A _2689_/B vssd1 vssd1 vccd1 vccd1 _2690_/A sky130_fd_sc_hd__and2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3104_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1991_ _2623_/B _1991_/B _2623_/D _1991_/D vssd1 vssd1 vccd1 vccd1 _2471_/D sky130_fd_sc_hd__or4_4
XFILLER_60_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2612_ _3150_/Q _2606_/X _2611_/X _3149_/Q vssd1 vssd1 vccd1 vccd1 _2612_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_62_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2543_ _2498_/X _2541_/X _2542_/X _2517_/X vssd1 vssd1 vccd1 vccd1 _3129_/D sky130_fd_sc_hd__o211a_1
X_2474_ _2474_/A _2474_/B vssd1 vssd1 vccd1 vccd1 _2547_/A sky130_fd_sc_hd__nor2_1
XFILLER_68_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3026_ _3028_/CLK _3026_/D vssd1 vssd1 vccd1 vccd1 _3026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2190_ _3035_/Q _2189_/X _2167_/X _3034_/Q vssd1 vssd1 vccd1 vccd1 _2190_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1974_ _3249_/Q vssd1 vssd1 vccd1 vccd1 _2457_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2526_ _2526_/A _2526_/B vssd1 vssd1 vccd1 vccd1 _2526_/Y sky130_fd_sc_hd__nand2_2
X_2457_ _2457_/A vssd1 vssd1 vccd1 vccd1 _2621_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2388_ _2096_/X _2387_/Y _2381_/X vssd1 vssd1 vccd1 vccd1 _3089_/D sky130_fd_sc_hd__a21oi_1
XFILLER_71_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3009_ _3100_/CLK _3009_/D vssd1 vssd1 vccd1 vccd1 _3009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1690_ _3416_/A _2929_/C _2867_/A vssd1 vssd1 vccd1 vccd1 _3247_/D sky130_fd_sc_hd__a21oi_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _2351_/A vssd1 vssd1 vccd1 vccd1 _2311_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ _2239_/X _2240_/Y _2241_/X vssd1 vssd1 vccd1 vccd1 _3044_/D sky130_fd_sc_hd__a21oi_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2173_ _2171_/Y _2172_/Y _2155_/X vssd1 vssd1 vccd1 vccd1 _3032_/D sky130_fd_sc_hd__a21oi_1
XFILLER_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1957_ _3004_/Q _1919_/X _1929_/X _3003_/Q vssd1 vssd1 vccd1 vccd1 _1957_/Y sky130_fd_sc_hd__a22oi_1
X_1888_ _3252_/Q _1888_/B _1888_/C _1836_/A vssd1 vssd1 vccd1 vccd1 _2267_/B sky130_fd_sc_hd__nor4b_1
X_2509_ _3124_/Q _2507_/X _2483_/X _3123_/Q _2939_/B vssd1 vssd1 vccd1 vccd1 _2509_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_14 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_471 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2860_ _3221_/Q _2853_/X _2859_/X _3220_/Q vssd1 vssd1 vccd1 vccd1 _2860_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1811_ _2742_/B _2905_/B vssd1 vssd1 vccd1 vccd1 _1811_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2791_ _2773_/X _2789_/X _2790_/X _2708_/X vssd1 vssd1 vccd1 vccd1 _3199_/D sky130_fd_sc_hd__o211a_1
X_1742_ _1804_/A vssd1 vssd1 vccd1 vccd1 _1960_/B sky130_fd_sc_hd__clkbuf_2
X_1673_ _2867_/A vssd1 vssd1 vccd1 vccd1 _1681_/A sky130_fd_sc_hd__clkbuf_2
X_3412_ _3412_/A _1666_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _2500_/A vssd1 vssd1 vccd1 vccd1 _2526_/A sky130_fd_sc_hd__buf_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2156_ _2153_/Y _2154_/Y _2155_/X vssd1 vssd1 vccd1 vccd1 _3029_/D sky130_fd_sc_hd__a21oi_1
XFILLER_26_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2087_ _2085_/B _1878_/A _1823_/A _1949_/B _2128_/A vssd1 vssd1 vccd1 vccd1 _2248_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2989_ _3113_/CLK _2989_/D vssd1 vssd1 vccd1 vccd1 _3406_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2010_ _3008_/Q _1986_/X _1994_/X _3007_/Q vssd1 vssd1 vccd1 vccd1 _2010_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_82_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3269_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2912_ _2912_/A _2912_/B _2912_/C _2912_/D vssd1 vssd1 vccd1 vccd1 _2912_/X sky130_fd_sc_hd__or4_1
X_2843_ _2843_/A vssd1 vssd1 vccd1 vccd1 _2843_/X sky130_fd_sc_hd__clkbuf_2
X_2774_ _1829_/X _1739_/Y _2170_/D _2686_/A vssd1 vssd1 vccd1 vccd1 _2774_/X sky130_fd_sc_hd__a211o_1
X_1725_ _3255_/Q vssd1 vssd1 vccd1 vccd1 _1946_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1656_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1656_/Y sky130_fd_sc_hd__inv_2
X_1587_ _1587_/A vssd1 vssd1 vccd1 vccd1 _1587_/Y sky130_fd_sc_hd__inv_2
X_3363__5 vssd1 vssd1 vccd1 vccd1 _3363__5/HI _3363_/A sky130_fd_sc_hd__conb_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_316 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3257_ _3270_/CLK _3257_/D vssd1 vssd1 vccd1 vccd1 _3257_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _3038_/Q _2189_/X _2195_/X _3037_/Q vssd1 vssd1 vccd1 vccd1 _2208_/Y sky130_fd_sc_hd__a22oi_1
X_3188_ _3269_/CLK _3188_/D vssd1 vssd1 vccd1 vccd1 _3188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2139_ _2227_/A vssd1 vssd1 vccd1 vccd1 _2139_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2490_ _2508_/A vssd1 vssd1 vccd1 vccd1 _2524_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3111_ _3116_/CLK _3111_/D vssd1 vssd1 vccd1 vccd1 _3111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3042_ _3069_/CLK _3042_/D vssd1 vssd1 vccd1 vccd1 _3042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2826_ _2826_/A _3209_/Q vssd1 vssd1 vccd1 vccd1 _2826_/X sky130_fd_sc_hd__or2_1
X_2757_ _2754_/X _2756_/X _2638_/A vssd1 vssd1 vccd1 vccd1 _2757_/X sky130_fd_sc_hd__a21o_1
X_1708_ _2947_/A _3405_/A vssd1 vssd1 vccd1 vccd1 _1708_/X sky130_fd_sc_hd__or2_1
X_2688_ _3173_/Q _2687_/X _2483_/A _3172_/Q _2508_/A vssd1 vssd1 vccd1 vccd1 _2689_/B
+ sky130_fd_sc_hd__o221a_1
X_1639_ _1642_/A vssd1 vssd1 vccd1 vccd1 _1639_/Y sky130_fd_sc_hd__inv_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_14 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1990_ _2474_/B _1843_/B _2268_/B vssd1 vssd1 vccd1 vccd1 _1991_/D sky130_fd_sc_hd__a21oi_2
X_2611_ _2783_/A vssd1 vssd1 vccd1 vccd1 _2611_/X sky130_fd_sc_hd__clkbuf_2
X_2542_ _3129_/Q _2542_/B vssd1 vssd1 vccd1 vccd1 _2542_/X sky130_fd_sc_hd__or2_1
XFILLER_55_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2473_ _2471_/X _2472_/Y _2458_/X vssd1 vssd1 vccd1 vccd1 _3119_/D sky130_fd_sc_hd__a21oi_1
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3025_ _3028_/CLK _3025_/D vssd1 vssd1 vccd1 vccd1 _3025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2809_ _2175_/X _2808_/Y _2794_/X vssd1 vssd1 vccd1 vccd1 _3204_/D sky130_fd_sc_hd__a21oi_1
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_447 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1973_ _3005_/Q _1919_/X _1929_/X _3004_/Q vssd1 vssd1 vccd1 vccd1 _1973_/Y sky130_fd_sc_hd__a22oi_1
X_2525_ _2525_/A vssd1 vssd1 vccd1 vccd1 _3126_/D sky130_fd_sc_hd__clkbuf_1
X_2456_ _3115_/Q _2446_/X _2449_/X _3114_/Q vssd1 vssd1 vccd1 vccd1 _2456_/Y sky130_fd_sc_hd__a22oi_1
X_2387_ _3089_/Q _2383_/X _2386_/X _3088_/Q vssd1 vssd1 vccd1 vccd1 _2387_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_71_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3008_ _3104_/CLK _3008_/D vssd1 vssd1 vccd1 vccd1 _3008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_73 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ _2256_/Y _2307_/Y _2309_/X vssd1 vssd1 vccd1 vccd1 _3061_/D sky130_fd_sc_hd__a21oi_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _2294_/A vssd1 vssd1 vccd1 vccd1 _2241_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2172_ _3032_/Q _2159_/X _2167_/X _3031_/Q vssd1 vssd1 vccd1 vccd1 _2172_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1956_ _1956_/A vssd1 vssd1 vccd1 vccd1 _1956_/X sky130_fd_sc_hd__buf_2
XFILLER_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1887_ _1940_/A _1887_/B vssd1 vssd1 vccd1 vccd1 _2693_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2508_ _2508_/A vssd1 vssd1 vccd1 vccd1 _2939_/B sky130_fd_sc_hd__clkbuf_2
X_2439_ _1905_/Y _2438_/Y _2430_/X vssd1 vssd1 vccd1 vccd1 _3108_/D sky130_fd_sc_hd__a21oi_1
XFILLER_56_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1810_ _1896_/A vssd1 vssd1 vccd1 vccd1 _2905_/B sky130_fd_sc_hd__clkbuf_2
X_2790_ _3199_/Q _2842_/B vssd1 vssd1 vccd1 vccd1 _2790_/X sky130_fd_sc_hd__or2_1
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1741_ _1825_/B vssd1 vssd1 vccd1 vccd1 _1960_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_362 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1672_ _2980_/Q _1672_/B vssd1 vssd1 vccd1 vccd1 _2980_/D sky130_fd_sc_hd__nor2_1
X_3411_ _3411_/A _1665_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _2677_/B _2474_/A _2710_/A _2223_/Y _2547_/C vssd1 vssd1 vccd1 vccd1 _2224_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _2155_/A vssd1 vssd1 vccd1 vccd1 _2155_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2086_ _2086_/A vssd1 vssd1 vccd1 vccd1 _2128_/A sky130_fd_sc_hd__buf_2
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3444__70 vssd1 vssd1 vccd1 vccd1 _3444__70/HI _3444_/A sky130_fd_sc_hd__conb_1
X_2988_ _3253_/CLK _2988_/D vssd1 vssd1 vccd1 vccd1 _3405_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1939_ _2537_/B _2537_/C vssd1 vssd1 vccd1 vccd1 _1939_/Y sky130_fd_sc_hd__nand2_1
X_3372__14 vssd1 vssd1 vccd1 vccd1 _3372__14/HI _3372_/A sky130_fd_sc_hd__conb_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2911_ _2472_/B _2909_/X _2910_/X _2843_/X vssd1 vssd1 vccd1 vccd1 _3240_/D sky130_fd_sc_hd__o211a_1
X_2842_ _3215_/Q _2842_/B vssd1 vssd1 vccd1 vccd1 _2842_/X sky130_fd_sc_hd__or2_1
X_2773_ _2773_/A vssd1 vssd1 vccd1 vccd1 _2773_/X sky130_fd_sc_hd__clkbuf_2
X_1724_ _1924_/B _1924_/A vssd1 vssd1 vccd1 vccd1 _1879_/A sky130_fd_sc_hd__and2b_1
X_1655_ _1661_/A vssd1 vssd1 vccd1 vccd1 _1660_/A sky130_fd_sc_hd__buf_2
X_1586_ _1587_/A vssd1 vssd1 vccd1 vccd1 _1586_/Y sky130_fd_sc_hd__inv_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3270_/CLK _3256_/D vssd1 vssd1 vccd1 vccd1 _3256_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _2835_/A _2477_/A _2205_/Y _2206_/X _1898_/X vssd1 vssd1 vccd1 vccd1 _2207_/Y
+ sky130_fd_sc_hd__o41ai_4
X_3187_ _3269_/CLK _3187_/D vssd1 vssd1 vccd1 vccd1 _3187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2138_ _2492_/C _2619_/C _2028_/X vssd1 vssd1 vccd1 vccd1 _2138_/Y sky130_fd_sc_hd__o21ai_1
X_2069_ _1880_/X _2122_/B _2681_/A _1829_/X vssd1 vssd1 vccd1 vccd1 _2915_/B sky130_fd_sc_hd__a22o_1
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3110_ _3116_/CLK _3110_/D vssd1 vssd1 vccd1 vccd1 _3110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3041_ _3069_/CLK _3041_/D vssd1 vssd1 vccd1 vccd1 _3041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2825_ _2825_/A _2825_/B _2885_/B _2901_/C vssd1 vssd1 vccd1 vccd1 _2825_/X sky130_fd_sc_hd__or4_1
X_2756_ _2756_/A _2756_/B _2756_/C _2901_/C vssd1 vssd1 vccd1 vccd1 _2756_/X sky130_fd_sc_hd__or4_1
X_1707_ _2962_/A vssd1 vssd1 vccd1 vccd1 _2947_/A sky130_fd_sc_hd__clkbuf_2
X_2687_ _2687_/A vssd1 vssd1 vccd1 vccd1 _2687_/X sky130_fd_sc_hd__clkbuf_2
X_1638_ _1642_/A vssd1 vssd1 vccd1 vccd1 _1638_/Y sky130_fd_sc_hd__inv_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ _1575_/A vssd1 vssd1 vccd1 vccd1 _1574_/A sky130_fd_sc_hd__buf_6
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _3244_/CLK _3239_/D vssd1 vssd1 vccd1 vccd1 _3239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_438 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2610_ _1819_/X _2492_/B _2693_/D _2609_/X vssd1 vssd1 vccd1 vccd1 _3149_/D sky130_fd_sc_hd__o31a_1
X_2541_ _1997_/Y _2539_/X _2540_/X _3128_/Q vssd1 vssd1 vccd1 vccd1 _2541_/X sky130_fd_sc_hd__o2bb2a_1
X_2472_ _3119_/Q _2472_/B vssd1 vssd1 vccd1 vccd1 _2472_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3024_ _3028_/CLK _3024_/D vssd1 vssd1 vccd1 vccd1 _3024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3194_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2808_ _3204_/Q _2804_/X _2807_/X _3203_/Q vssd1 vssd1 vccd1 vccd1 _2808_/Y sky130_fd_sc_hd__a22oi_1
X_2739_ _3187_/Q _2520_/X _2522_/X _3186_/Q vssd1 vssd1 vccd1 vccd1 _2740_/C sky130_fd_sc_hd__o22a_1
XFILLER_3_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1972_ _1962_/X _1971_/X _1861_/X vssd1 vssd1 vccd1 vccd1 _1972_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_60_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2524_ _2524_/A _2524_/B _2524_/C vssd1 vssd1 vccd1 vccd1 _2525_/A sky130_fd_sc_hd__and3_1
X_2455_ _1839_/Y _2454_/Y _2443_/X vssd1 vssd1 vccd1 vccd1 _3114_/D sky130_fd_sc_hd__a21oi_1
X_2386_ _2406_/A vssd1 vssd1 vccd1 vccd1 _2386_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3007_ _3104_/CLK _3007_/D vssd1 vssd1 vccd1 vccd1 _3007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3378__20 vssd1 vssd1 vccd1 vccd1 _3378__20/HI _3378_/A sky130_fd_sc_hd__conb_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _3044_/Q _2218_/X _2227_/X _3043_/Q vssd1 vssd1 vccd1 vccd1 _2240_/Y sky130_fd_sc_hd__a22oi_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2171_ _1934_/Y _2584_/D _2028_/X vssd1 vssd1 vccd1 vccd1 _2171_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1955_ _2738_/A _2471_/B _2471_/C _1954_/X vssd1 vssd1 vccd1 vccd1 _1956_/A sky130_fd_sc_hd__or4b_1
X_1886_ _2061_/D vssd1 vssd1 vccd1 vccd1 _1940_/A sky130_fd_sc_hd__clkbuf_2
X_2507_ _2761_/A vssd1 vssd1 vccd1 vccd1 _2507_/X sky130_fd_sc_hd__clkbuf_2
X_2438_ _3108_/Q _2432_/X _2435_/X _3107_/Q vssd1 vssd1 vccd1 vccd1 _2438_/Y sky130_fd_sc_hd__a22oi_1
X_2369_ _3083_/Q _2365_/X _2368_/X _3082_/Q vssd1 vssd1 vccd1 vccd1 _2369_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_56_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_470 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1740_ _1909_/A vssd1 vssd1 vccd1 vccd1 _2061_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1671_ _2867_/A vssd1 vssd1 vccd1 vccd1 _1672_/B sky130_fd_sc_hd__buf_2
X_3410_ _3410_/A _1664_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2223_ _2223_/A _2223_/B vssd1 vssd1 vccd1 vccd1 _2223_/Y sky130_fd_sc_hd__nor2_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _3029_/Q _2132_/X _2139_/X _3028_/Q vssd1 vssd1 vccd1 vccd1 _2154_/Y sky130_fd_sc_hd__a22oi_1
X_2085_ _2085_/A _2085_/B _2262_/B vssd1 vssd1 vccd1 vccd1 _2248_/A sky130_fd_sc_hd__or3_1
XFILLER_53_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2987_ _3152_/CLK _2987_/D vssd1 vssd1 vccd1 vccd1 _2987_/Q sky130_fd_sc_hd__dfxtp_1
X_1938_ _1835_/C _2122_/B _2681_/A _2583_/A vssd1 vssd1 vccd1 vccd1 _2467_/A sky130_fd_sc_hd__a22o_2
X_1869_ _1946_/A _1893_/B _1913_/B vssd1 vssd1 vccd1 vccd1 _2178_/A sky130_fd_sc_hd__nand3b_2
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2910_ _3240_/Q _2924_/B vssd1 vssd1 vccd1 vccd1 _2910_/X sky130_fd_sc_hd__or2_1
X_2841_ _2540_/X _3214_/Q _2274_/X _2819_/D vssd1 vssd1 vccd1 vccd1 _2841_/X sky130_fd_sc_hd__o22a_1
XFILLER_78_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2772_ _2080_/X _2771_/X _2394_/X vssd1 vssd1 vccd1 vccd1 _3194_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3113_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1723_ _3252_/Q vssd1 vssd1 vccd1 vccd1 _1924_/A sky130_fd_sc_hd__clkbuf_1
X_1654_ _1654_/A vssd1 vssd1 vccd1 vccd1 _1654_/Y sky130_fd_sc_hd__inv_2
X_1585_ _1587_/A vssd1 vssd1 vccd1 vccd1 _1585_/Y sky130_fd_sc_hd__inv_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3255_/CLK _3255_/D vssd1 vssd1 vccd1 vccd1 _3255_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2206_ _1999_/A _2223_/B _2199_/B _2116_/B _2005_/Y vssd1 vssd1 vccd1 vccd1 _2206_/X
+ sky130_fd_sc_hd__a311o_1
X_3186_ _3269_/CLK _3186_/D vssd1 vssd1 vccd1 vccd1 _3186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2137_ _2137_/A _2728_/B vssd1 vssd1 vccd1 vccd1 _2619_/C sky130_fd_sc_hd__nand2_2
XFILLER_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_384 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2068_ _2079_/B vssd1 vssd1 vccd1 vccd1 _2211_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3040_ _3069_/CLK _3040_/D vssd1 vssd1 vccd1 vccd1 _3040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2824_ _2810_/Y _2823_/Y _2817_/X vssd1 vssd1 vccd1 vccd1 _3209_/D sky130_fd_sc_hd__a21oi_1
X_2755_ _2472_/B _2753_/X _2754_/X _2699_/C _2722_/X vssd1 vssd1 vccd1 vccd1 _3190_/D
+ sky130_fd_sc_hd__o221a_1
X_1706_ _1696_/X _3405_/A _1700_/X _1705_/X vssd1 vssd1 vccd1 vccd1 _2987_/D sky130_fd_sc_hd__o211a_1
X_2686_ _2686_/A _2686_/B _2686_/C _2137_/A vssd1 vssd1 vccd1 vccd1 _2689_/A sky130_fd_sc_hd__or4b_1
X_1637_ _1637_/A vssd1 vssd1 vccd1 vccd1 _1642_/A sky130_fd_sc_hd__buf_4
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ _1568_/A vssd1 vssd1 vccd1 vccd1 _1568_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _3241_/CLK _3238_/D vssd1 vssd1 vccd1 vccd1 _3238_/Q sky130_fd_sc_hd__dfxtp_1
X_3169_ _3185_/CLK _3169_/D vssd1 vssd1 vccd1 vccd1 _3169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2540_ _2941_/S vssd1 vssd1 vccd1 vccd1 _2540_/X sky130_fd_sc_hd__buf_2
XFILLER_5_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2471_ _2848_/A _2471_/B _2471_/C _2471_/D vssd1 vssd1 vccd1 vccd1 _2471_/X sky130_fd_sc_hd__or4_4
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3023_ _3028_/CLK _3023_/D vssd1 vssd1 vccd1 vccd1 _3023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3402__44 vssd1 vssd1 vccd1 vccd1 _3402__44/HI _3402_/A sky130_fd_sc_hd__conb_1
X_2807_ _2874_/A vssd1 vssd1 vccd1 vccd1 _2807_/X sky130_fd_sc_hd__clkbuf_2
X_2738_ _2738_/A _2912_/D _2738_/C _2738_/D vssd1 vssd1 vccd1 vccd1 _2740_/B sky130_fd_sc_hd__or4_1
X_2669_ _2769_/A _2669_/B _2669_/C vssd1 vssd1 vccd1 vccd1 _2670_/A sky130_fd_sc_hd__and3_1
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_61 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1971_ _2677_/B _2474_/A _2710_/A _2912_/A _2623_/C vssd1 vssd1 vccd1 vccd1 _1971_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2523_ _3126_/Q _2520_/X _2522_/X _3125_/Q vssd1 vssd1 vccd1 vccd1 _2524_/C sky130_fd_sc_hd__o22a_1
X_2454_ _3114_/Q _2446_/X _2449_/X _3113_/Q vssd1 vssd1 vccd1 vccd1 _2454_/Y sky130_fd_sc_hd__a22oi_1
X_2385_ _2100_/Y _2384_/Y _2381_/X vssd1 vssd1 vccd1 vccd1 _3088_/D sky130_fd_sc_hd__a21oi_1
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3006_ _3104_/CLK _3006_/D vssd1 vssd1 vccd1 vccd1 _3006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_228 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3465__91 vssd1 vssd1 vccd1 vccd1 _3465__91/HI _3465_/A sky130_fd_sc_hd__conb_1
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_73 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3393__35 vssd1 vssd1 vccd1 vccd1 _3393__35/HI _3393_/A sky130_fd_sc_hd__conb_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_438 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2170_ _2170_/A _2681_/B _2170_/C _2170_/D vssd1 vssd1 vccd1 vccd1 _2584_/D sky130_fd_sc_hd__or4_4
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1954_ _1981_/A _2129_/B _1953_/X _1903_/A vssd1 vssd1 vccd1 vccd1 _1954_/X sky130_fd_sc_hd__o211a_1
X_1885_ _1879_/A _1968_/A _1880_/X _1963_/A vssd1 vssd1 vccd1 vccd1 _2756_/B sky130_fd_sc_hd__a22o_1
X_2506_ _2748_/A _2199_/B _2274_/B _1934_/Y _2552_/C vssd1 vssd1 vccd1 vccd1 _2506_/X
+ sky130_fd_sc_hd__a2111o_1
X_2437_ _1916_/X _2436_/Y _2430_/X vssd1 vssd1 vccd1 vccd1 _3107_/D sky130_fd_sc_hd__a21oi_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2368_ _2406_/A vssd1 vssd1 vccd1 vccd1 _2368_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2299_ _2276_/Y _2298_/Y _2294_/X vssd1 vssd1 vccd1 vccd1 _3057_/D sky130_fd_sc_hd__a21oi_1
XFILLER_56_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1670_ _3249_/Q vssd1 vssd1 vccd1 vccd1 _2867_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _2046_/A _2623_/C _2477_/A _2885_/B vssd1 vssd1 vccd1 vccd1 _2222_/X sky130_fd_sc_hd__a211o_1
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2153_ _2835_/A _2532_/A _1916_/D _1992_/X vssd1 vssd1 vccd1 vccd1 _2153_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_19_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2084_ _2901_/A _2567_/C vssd1 vssd1 vccd1 vccd1 _2734_/C sky130_fd_sc_hd__or2_1
XFILLER_34_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2986_ _3248_/CLK _2986_/D vssd1 vssd1 vccd1 vccd1 _3416_/A sky130_fd_sc_hd__dfxtp_1
X_1937_ _1937_/A vssd1 vssd1 vccd1 vccd1 _2583_/A sky130_fd_sc_hd__clkbuf_2
X_1868_ _1868_/A vssd1 vssd1 vccd1 vccd1 _2268_/A sky130_fd_sc_hd__clkbuf_2
X_1799_ _1913_/B _1953_/D _1913_/C vssd1 vssd1 vccd1 vccd1 _2001_/A sky130_fd_sc_hd__nor3_2
X_3469_ _3469_/A _1648_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
XFILLER_67_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3013_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3435__61 vssd1 vssd1 vccd1 vccd1 _3435__61/HI _3435_/A sky130_fd_sc_hd__conb_1
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2840_ _2207_/Y _2839_/Y _2817_/X vssd1 vssd1 vccd1 vccd1 _3214_/D sky130_fd_sc_hd__a21oi_1
XFILLER_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2771_ _3194_/Q _2497_/A _2290_/X _3193_/Q vssd1 vssd1 vccd1 vccd1 _2771_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1722_ _3251_/Q vssd1 vssd1 vccd1 vccd1 _1924_/B sky130_fd_sc_hd__clkbuf_1
X_1653_ _1654_/A vssd1 vssd1 vccd1 vccd1 _1653_/Y sky130_fd_sc_hd__inv_2
X_1584_ _1587_/A vssd1 vssd1 vccd1 vccd1 _1584_/Y sky130_fd_sc_hd__inv_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _3255_/CLK _3254_/D vssd1 vssd1 vccd1 vccd1 _3254_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2205_/A _2731_/A vssd1 vssd1 vccd1 vccd1 _2205_/Y sky130_fd_sc_hd__nand2_1
X_3185_ _3185_/CLK _3185_/D vssd1 vssd1 vccd1 vccd1 _3185_/Q sky130_fd_sc_hd__dfxtp_1
X_2136_ _2742_/A _2905_/C _2181_/B vssd1 vssd1 vccd1 vccd1 _2492_/C sky130_fd_sc_hd__or3_1
XFILLER_66_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2067_ _2067_/A vssd1 vssd1 vccd1 vccd1 _2819_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2969_ _2971_/A _3267_/Q vssd1 vssd1 vccd1 vccd1 _2969_/X sky130_fd_sc_hd__or2_1
XFILLER_1_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2823_ _3209_/Q _2804_/X _2807_/X _3208_/Q vssd1 vssd1 vccd1 vccd1 _2823_/Y sky130_fd_sc_hd__a22oi_1
X_2754_ _2826_/A _3190_/Q vssd1 vssd1 vccd1 vccd1 _2754_/X sky130_fd_sc_hd__or2_1
X_1705_ _1705_/A _2987_/Q vssd1 vssd1 vccd1 vccd1 _1705_/X sky130_fd_sc_hd__or2_1
X_2685_ _2638_/X _2682_/X _2684_/X _2632_/X vssd1 vssd1 vccd1 vccd1 _3172_/D sky130_fd_sc_hd__o211a_1
X_1636_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1636_/Y sky130_fd_sc_hd__inv_2
X_1567_ _1568_/A vssd1 vssd1 vccd1 vccd1 _1567_/Y sky130_fd_sc_hd__inv_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3241_/CLK _3237_/D vssd1 vssd1 vccd1 vccd1 _3237_/Q sky130_fd_sc_hd__dfxtp_1
X_3168_ _3168_/CLK _3168_/D vssd1 vssd1 vccd1 vccd1 _3168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2119_ _1838_/A _1804_/X _2116_/Y _2118_/X _1812_/X vssd1 vssd1 vccd1 vccd1 _2119_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3099_ _3103_/CLK _3099_/D vssd1 vssd1 vccd1 vccd1 _3099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_196 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2470_ _2738_/A vssd1 vssd1 vccd1 vccd1 _2848_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3022_ _3082_/CLK _3022_/D vssd1 vssd1 vccd1 vccd1 _3022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_358 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3399__41 vssd1 vssd1 vccd1 vccd1 _3399__41/HI _3399_/A sky130_fd_sc_hd__conb_1
X_2806_ _2803_/Y _2805_/Y _2794_/X vssd1 vssd1 vccd1 vccd1 _3203_/D sky130_fd_sc_hd__a21oi_1
X_2737_ _2737_/A vssd1 vssd1 vccd1 vccd1 _3186_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3241_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2668_ _3168_/Q _2520_/X _2522_/X _3167_/Q vssd1 vssd1 vccd1 vccd1 _2669_/C sky130_fd_sc_hd__o22a_1
X_1619_ _1637_/A vssd1 vssd1 vccd1 vccd1 _1624_/A sky130_fd_sc_hd__clkbuf_4
X_2599_ _3145_/Q _2580_/X _2586_/X _3144_/Q vssd1 vssd1 vccd1 vccd1 _2599_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_59_425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_344 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1970_ _2198_/A vssd1 vssd1 vccd1 vccd1 _2912_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2522_ _2767_/A vssd1 vssd1 vccd1 vccd1 _2522_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2453_ _2801_/B _2452_/Y _2443_/X vssd1 vssd1 vccd1 vccd1 _3113_/D sky130_fd_sc_hd__a21oi_1
X_2384_ _3088_/Q _2383_/X _2368_/X _3087_/Q vssd1 vssd1 vccd1 vccd1 _2384_/Y sky130_fd_sc_hd__a22oi_1
Xinput2 la1_data_in[0] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3005_ _3104_/CLK _3005_/D vssd1 vssd1 vccd1 vccd1 _3005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1953_ _2034_/D _1953_/B _1960_/B _1953_/D vssd1 vssd1 vccd1 vccd1 _1953_/X sky130_fd_sc_hd__or4_1
X_3369__11 vssd1 vssd1 vccd1 vccd1 _3369__11/HI _3369_/A sky130_fd_sc_hd__conb_1
X_1884_ _1882_/X _1883_/Y _1853_/X vssd1 vssd1 vccd1 vccd1 _2998_/D sky130_fd_sc_hd__a21oi_1
X_3366__8 vssd1 vssd1 vccd1 vccd1 _3366__8/HI _3366_/A sky130_fd_sc_hd__conb_1
X_2505_ _2498_/X _2501_/X _2504_/X _2394_/X vssd1 vssd1 vccd1 vccd1 _3123_/D sky130_fd_sc_hd__o211a_1
X_2436_ _3107_/Q _2432_/X _2435_/X _3106_/Q vssd1 vssd1 vccd1 vccd1 _2436_/Y sky130_fd_sc_hd__a22oi_1
X_2367_ _2138_/Y _2366_/Y _2362_/X vssd1 vssd1 vccd1 vccd1 _3082_/D sky130_fd_sc_hd__a21oi_1
XFILLER_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2298_ _3057_/Q _2297_/X _2277_/X _3056_/Q vssd1 vssd1 vccd1 vccd1 _2298_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_64_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3270_ _3270_/CLK _3270_/D vssd1 vssd1 vccd1 vccd1 _3409_/A sky130_fd_sc_hd__dfxtp_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _1940_/A _2122_/B _1997_/B vssd1 vssd1 vccd1 vccd1 _2885_/B sky130_fd_sc_hd__a21o_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2152_ _2152_/A vssd1 vssd1 vccd1 vccd1 _2532_/A sky130_fd_sc_hd__buf_2
X_2083_ _2080_/X _2082_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _3017_/D sky130_fd_sc_hd__o21a_1
XFILLER_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2985_ _3248_/CLK _2985_/D vssd1 vssd1 vccd1 vccd1 _3415_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1936_ _1936_/A vssd1 vssd1 vccd1 vccd1 _1937_/A sky130_fd_sc_hd__inv_2
X_1867_ _2012_/A _2477_/C vssd1 vssd1 vccd1 vccd1 _2686_/C sky130_fd_sc_hd__or2_1
X_1798_ _1806_/D vssd1 vssd1 vccd1 vccd1 _1913_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3468_ _3468_/A _1647_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
X_3399_ _3399_/A _1602_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_76_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2419_ _3101_/Q _2418_/X _2406_/X _3100_/Q vssd1 vssd1 vccd1 vccd1 _2419_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_72_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3450__76 vssd1 vssd1 vccd1 vccd1 _3450__76/HI _3450_/A sky130_fd_sc_hd__conb_1
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2770_ _2770_/A vssd1 vssd1 vccd1 vccd1 _3193_/D sky130_fd_sc_hd__clkbuf_1
X_1721_ _1998_/A _1909_/A _1825_/B vssd1 vssd1 vccd1 vccd1 _1963_/A sky130_fd_sc_hd__nor3b_2
XFILLER_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1652_ _1654_/A vssd1 vssd1 vccd1 vccd1 _1652_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1583_ _1587_/A vssd1 vssd1 vccd1 vccd1 _1583_/Y sky130_fd_sc_hd__inv_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3253_/CLK _3253_/D vssd1 vssd1 vccd1 vccd1 _3253_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _3242_/CLK _3184_/D vssd1 vssd1 vccd1 vccd1 _3184_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _2204_/A vssd1 vssd1 vccd1 vccd1 _2477_/A sky130_fd_sc_hd__clkbuf_4
X_2135_ _2094_/B _1910_/A _1807_/A _1937_/A _1961_/A vssd1 vssd1 vccd1 vccd1 _2181_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_66_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2066_ _2064_/X _2065_/Y _2043_/X vssd1 vssd1 vccd1 vccd1 _3014_/D sky130_fd_sc_hd__a21oi_1
XFILLER_22_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2968_ _1696_/A _3267_/Q _2959_/X _2967_/X vssd1 vssd1 vccd1 vccd1 _3266_/D sky130_fd_sc_hd__o211a_1
X_1919_ _2132_/A vssd1 vssd1 vccd1 vccd1 _1919_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2899_ _3237_/Q _2542_/B _2712_/X _3236_/Q _2713_/X vssd1 vssd1 vccd1 vccd1 _2899_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_14 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_386 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2822_ _2822_/A vssd1 vssd1 vccd1 vccd1 _3208_/D sky130_fd_sc_hd__clkbuf_1
X_2753_ _2157_/B _2915_/B _2752_/Y _3189_/Q _2540_/X vssd1 vssd1 vccd1 vccd1 _2753_/X
+ sky130_fd_sc_hd__o32a_1
X_1704_ _2962_/A vssd1 vssd1 vccd1 vccd1 _1705_/A sky130_fd_sc_hd__buf_2
X_2684_ _3172_/Q _2842_/B vssd1 vssd1 vccd1 vccd1 _2684_/X sky130_fd_sc_hd__or2_1
X_1635_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1635_/Y sky130_fd_sc_hd__inv_2
X_1566_ _1568_/A vssd1 vssd1 vccd1 vccd1 _1566_/Y sky130_fd_sc_hd__inv_2
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3236_ _3241_/CLK _3236_/D vssd1 vssd1 vccd1 vccd1 _3236_/Q sky130_fd_sc_hd__dfxtp_1
X_3167_ _3270_/CLK _3167_/D vssd1 vssd1 vccd1 vccd1 _3167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3098_ _3100_/CLK _3098_/D vssd1 vssd1 vccd1 vccd1 _3098_/Q sky130_fd_sc_hd__dfxtp_1
X_2118_ _2825_/B _2231_/B vssd1 vssd1 vccd1 vccd1 _2118_/X sky130_fd_sc_hd__and2b_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2049_ _2045_/X _2046_/Y _2047_/X _2048_/X vssd1 vssd1 vccd1 vccd1 _2049_/X sky130_fd_sc_hd__a31o_1
XFILLER_80_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3420__46 vssd1 vssd1 vccd1 vccd1 _3420__46/HI _3420_/A sky130_fd_sc_hd__conb_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3021_ _3092_/CLK _3021_/D vssd1 vssd1 vccd1 vccd1 _3021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2805_ _3203_/Q _2804_/X _2783_/X _3202_/Q vssd1 vssd1 vccd1 vccd1 _2805_/Y sky130_fd_sc_hd__a22oi_1
X_2736_ _2736_/A _2736_/B vssd1 vssd1 vccd1 vccd1 _2737_/A sky130_fd_sc_hd__and2_1
X_2667_ _2667_/A _2912_/C _2667_/C _2667_/D vssd1 vssd1 vccd1 vccd1 _2669_/B sky130_fd_sc_hd__or4_1
X_1618_ _1618_/A vssd1 vssd1 vccd1 vccd1 _1618_/Y sky130_fd_sc_hd__inv_2
X_2598_ _1857_/A _2596_/Y _2597_/X vssd1 vssd1 vccd1 vccd1 _3144_/D sky130_fd_sc_hd__a21boi_1
X_1549_ _1549_/A vssd1 vssd1 vccd1 vccd1 _1549_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3219_ _3234_/CLK _3219_/D vssd1 vssd1 vccd1 vccd1 _3219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2521_ _2624_/A vssd1 vssd1 vccd1 vccd1 _2767_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2452_ _3113_/Q _2446_/X _2449_/X _3112_/Q vssd1 vssd1 vccd1 vccd1 _2452_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_5_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2383_ _2432_/A vssd1 vssd1 vccd1 vccd1 _2383_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3004_ _3104_/CLK _3004_/D vssd1 vssd1 vccd1 vccd1 _3004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2719_ _2212_/A _2474_/B _2716_/Y _2718_/Y _1681_/A vssd1 vssd1 vccd1 vccd1 _3180_/D
+ sky130_fd_sc_hd__a311oi_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3456__82 vssd1 vssd1 vccd1 vccd1 _3456__82/HI _3456_/A sky130_fd_sc_hd__conb_1
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1952_ _2003_/A _2012_/A _1980_/C vssd1 vssd1 vccd1 vccd1 _2471_/C sky130_fd_sc_hd__a21o_2
X_1883_ _2998_/Q _1863_/X _1874_/X _2997_/Q vssd1 vssd1 vccd1 vccd1 _1883_/Y sky130_fd_sc_hd__a22oi_1
X_3384__26 vssd1 vssd1 vccd1 vccd1 _3384__26/HI _3384_/A sky130_fd_sc_hd__conb_1
X_2504_ _3123_/Q _2542_/B vssd1 vssd1 vccd1 vccd1 _2504_/X sky130_fd_sc_hd__or2_1
X_2435_ _2559_/A vssd1 vssd1 vccd1 vccd1 _2435_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2366_ _3082_/Q _2365_/X _2354_/X _3081_/Q vssd1 vssd1 vccd1 vccd1 _2366_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2297_ _2351_/A vssd1 vssd1 vccd1 vccd1 _2297_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2217_/Y _2219_/Y _2214_/X vssd1 vssd1 vccd1 vccd1 _3040_/D sky130_fd_sc_hd__a21oi_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2151_ _2149_/Y _2150_/Y _2125_/X vssd1 vssd1 vccd1 vccd1 _3028_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2082_ _3017_/Q _2081_/X _2020_/X _3016_/Q vssd1 vssd1 vccd1 vccd1 _2082_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2984_ _3248_/CLK _2984_/D vssd1 vssd1 vccd1 vccd1 _3414_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1935_ _1935_/A vssd1 vssd1 vccd1 vccd1 _2681_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1866_ _1866_/A vssd1 vssd1 vccd1 vccd1 _2012_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1797_ _1888_/C vssd1 vssd1 vccd1 vccd1 _1913_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3467_ _3467_/A _1646_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
X_3398_ _3398_/A _1601_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
X_2418_ _2432_/A vssd1 vssd1 vccd1 vccd1 _2418_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2349_ _2362_/A vssd1 vssd1 vccd1 vccd1 _2349_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_336 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3426__52 vssd1 vssd1 vccd1 vccd1 _3426__52/HI _3426_/A sky130_fd_sc_hd__conb_1
XFILLER_43_262 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1720_ _3255_/Q vssd1 vssd1 vccd1 vccd1 _1825_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1651_ _1654_/A vssd1 vssd1 vccd1 vccd1 _1651_/Y sky130_fd_sc_hd__inv_2
X_1582_ _1606_/A vssd1 vssd1 vccd1 vccd1 _1587_/A sky130_fd_sc_hd__buf_4
XFILLER_3_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3255_/CLK _3252_/D vssd1 vssd1 vccd1 vccd1 _3252_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2203_ _2201_/X _2202_/Y _2185_/X vssd1 vssd1 vccd1 vccd1 _3037_/D sky130_fd_sc_hd__a21oi_1
X_3183_ _3248_/CLK _3183_/D vssd1 vssd1 vccd1 vccd1 _3183_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2134_ _2131_/Y _2133_/Y _2125_/X vssd1 vssd1 vccd1 vccd1 _3025_/D sky130_fd_sc_hd__a21oi_1
XFILLER_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2065_ _3014_/Q _2050_/X _2055_/X _3013_/Q vssd1 vssd1 vccd1 vccd1 _2065_/Y sky130_fd_sc_hd__a22oi_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3070_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2967_ _2971_/A _3266_/Q vssd1 vssd1 vccd1 vccd1 _2967_/X sky130_fd_sc_hd__or2_1
X_2898_ _2743_/C _2788_/X _2897_/X vssd1 vssd1 vccd1 vccd1 _3236_/D sky130_fd_sc_hd__o21a_1
X_1918_ _2296_/A vssd1 vssd1 vccd1 vccd1 _2132_/A sky130_fd_sc_hd__clkbuf_2
X_1849_ _2477_/C _2905_/C vssd1 vssd1 vccd1 vccd1 _1851_/B sky130_fd_sc_hd__or2_4
XFILLER_78_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2821_ _2907_/A _2821_/B _2821_/C vssd1 vssd1 vccd1 vccd1 _2822_/A sky130_fd_sc_hd__and3_1
XFILLER_76_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2752_ _2752_/A _2752_/B vssd1 vssd1 vccd1 vccd1 _2752_/Y sky130_fd_sc_hd__nand2_1
X_1703_ _2728_/A vssd1 vssd1 vccd1 vccd1 _2962_/A sky130_fd_sc_hd__clkbuf_2
X_2683_ _2683_/A vssd1 vssd1 vccd1 vccd1 _2842_/B sky130_fd_sc_hd__clkbuf_2
X_1634_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1634_/Y sky130_fd_sc_hd__inv_2
X_1565_ _1568_/A vssd1 vssd1 vccd1 vccd1 _1565_/Y sky130_fd_sc_hd__inv_2
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _3241_/CLK _3235_/D vssd1 vssd1 vccd1 vccd1 _3235_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _3270_/CLK _3166_/D vssd1 vssd1 vccd1 vccd1 _3166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2117_ _2537_/B _2262_/B _1823_/A _2747_/B _2198_/B vssd1 vssd1 vccd1 vccd1 _2231_/B
+ sky130_fd_sc_hd__o32a_1
X_3097_ _3100_/CLK _3097_/D vssd1 vssd1 vccd1 vccd1 _3097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2048_ _2765_/B vssd1 vssd1 vccd1 vccd1 _2048_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3020_ _3092_/CLK _3020_/D vssd1 vssd1 vccd1 vccd1 _3020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2804_ _2829_/A vssd1 vssd1 vccd1 vccd1 _2804_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2735_ _3186_/Q _2687_/X _2625_/A _3185_/Q _2393_/A vssd1 vssd1 vccd1 vccd1 _2736_/B
+ sky130_fd_sc_hd__o221a_1
X_2666_ _2467_/X _2664_/Y _2665_/X vssd1 vssd1 vccd1 vccd1 _3167_/D sky130_fd_sc_hd__a21oi_1
X_1617_ _1618_/A vssd1 vssd1 vccd1 vccd1 _1617_/Y sky130_fd_sc_hd__inv_2
X_2597_ _3144_/Q _2511_/A _2493_/X _3143_/Q _2929_/B vssd1 vssd1 vccd1 vccd1 _2597_/X
+ sky130_fd_sc_hd__o221a_1
X_1548_ _1549_/A vssd1 vssd1 vccd1 vccd1 _1548_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_31_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3168_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3218_ _3232_/CLK _3218_/D vssd1 vssd1 vccd1 vccd1 _3218_/Q sky130_fd_sc_hd__dfxtp_1
X_3149_ _3149_/CLK _3149_/D vssd1 vssd1 vccd1 vccd1 _3149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_316 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_419 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_474 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2520_ _2766_/A vssd1 vssd1 vccd1 vccd1 _2520_/X sky130_fd_sc_hd__clkbuf_2
X_2451_ _1862_/Y _2450_/Y _2443_/X vssd1 vssd1 vccd1 vccd1 _3112_/D sky130_fd_sc_hd__a21oi_1
XFILLER_5_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2382_ _2108_/X _2379_/Y _2381_/X vssd1 vssd1 vccd1 vccd1 _3087_/D sky130_fd_sc_hd__a21oi_1
XFILLER_49_460 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3003_ _3104_/CLK _3003_/D vssd1 vssd1 vccd1 vccd1 _3003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2718_ _3180_/Q _2924_/B _2493_/X _3179_/Q vssd1 vssd1 vccd1 vccd1 _2718_/Y sky130_fd_sc_hd__o22ai_1
X_2649_ _2846_/A vssd1 vssd1 vccd1 vccd1 _2649_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1951_ _1965_/A _1951_/B _2001_/A vssd1 vssd1 vccd1 vccd1 _1980_/C sky130_fd_sc_hd__and3_1
X_1882_ _2262_/B _2075_/A _2137_/A _2954_/A vssd1 vssd1 vccd1 vccd1 _1882_/X sky130_fd_sc_hd__a31o_1
X_2503_ _2761_/A vssd1 vssd1 vccd1 vccd1 _2542_/B sky130_fd_sc_hd__clkbuf_2
X_2434_ _1928_/Y _2433_/Y _2430_/X vssd1 vssd1 vccd1 vccd1 _3106_/D sky130_fd_sc_hd__a21oi_1
X_2365_ _2432_/A vssd1 vssd1 vccd1 vccd1 _2365_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2296_ _2296_/A vssd1 vssd1 vccd1 vccd1 _2351_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2150_ _3028_/Q _2132_/X _2139_/X _3027_/Q vssd1 vssd1 vccd1 vccd1 _2150_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2081_ _2871_/A vssd1 vssd1 vccd1 vccd1 _2081_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_400 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2983_ _3250_/CLK _2983_/D vssd1 vssd1 vccd1 vccd1 _3413_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1934_ _2085_/A _1856_/A _1887_/B vssd1 vssd1 vccd1 vccd1 _1934_/Y sky130_fd_sc_hd__o21ai_4
X_1865_ _1862_/Y _1864_/Y _1853_/X vssd1 vssd1 vccd1 vccd1 _2996_/D sky130_fd_sc_hd__a21oi_1
X_1796_ _1879_/A _2026_/B _1795_/X _1834_/A vssd1 vssd1 vccd1 vccd1 _2075_/A sky130_fd_sc_hd__o22a_2
X_3466_ _3466_/A _1645_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
X_2417_ _2009_/X _2415_/Y _2416_/X vssd1 vssd1 vccd1 vccd1 _3100_/D sky130_fd_sc_hd__a21oi_1
X_3397_ _3397_/A _1599_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_69_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2348_ _3076_/Q _2337_/X _2341_/X _3075_/Q vssd1 vssd1 vccd1 vccd1 _2348_/Y sky130_fd_sc_hd__a22oi_1
X_2279_ _2276_/Y _2278_/Y _2265_/X vssd1 vssd1 vccd1 vccd1 _3051_/D sky130_fd_sc_hd__a21oi_1
XFILLER_16_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_68 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3441__67 vssd1 vssd1 vccd1 vccd1 _3441__67/HI _3441_/A sky130_fd_sc_hd__conb_1
X_1650_ _1654_/A vssd1 vssd1 vccd1 vccd1 _1650_/Y sky130_fd_sc_hd__inv_2
X_1581_ input1/X vssd1 vssd1 vccd1 vccd1 _1606_/A sky130_fd_sc_hd__clkbuf_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3253_/CLK _3251_/D vssd1 vssd1 vccd1 vccd1 _3251_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _3037_/Q _2189_/X _2195_/X _3036_/Q vssd1 vssd1 vccd1 vccd1 _2202_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3182_ _3248_/CLK _3182_/D vssd1 vssd1 vccd1 vccd1 _3182_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2133_ _3025_/Q _2132_/X _2102_/X _3024_/Q vssd1 vssd1 vccd1 vccd1 _2133_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2064_ _2584_/A _2519_/C _2064_/C vssd1 vssd1 vccd1 vccd1 _2064_/X sky130_fd_sc_hd__or3_4
XFILLER_22_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2966_ _2954_/X _3266_/Q _2959_/X _2965_/X vssd1 vssd1 vccd1 vccd1 _3265_/D sky130_fd_sc_hd__o211a_1
X_2897_ _3236_/Q _2527_/X _2528_/X _3235_/Q _2524_/A vssd1 vssd1 vccd1 vccd1 _2897_/X
+ sky130_fd_sc_hd__o221a_1
X_1917_ _1917_/A vssd1 vssd1 vccd1 vccd1 _2296_/A sky130_fd_sc_hd__clkbuf_2
X_1848_ _1804_/X _1803_/A _1895_/A vssd1 vssd1 vccd1 vccd1 _2905_/C sky130_fd_sc_hd__a21oi_2
X_1779_ _2871_/A vssd1 vssd1 vccd1 vccd1 _2773_/A sky130_fd_sc_hd__buf_2
XFILLER_1_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3449_ _3449_/A _1618_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2820_ _3208_/Q _2766_/X _2767_/X _3207_/Q vssd1 vssd1 vccd1 vccd1 _2821_/C sky130_fd_sc_hd__o22a_1
X_2751_ _2751_/A vssd1 vssd1 vccd1 vccd1 _3189_/D sky130_fd_sc_hd__clkbuf_1
X_1702_ _2538_/A vssd1 vssd1 vccd1 vccd1 _2728_/A sky130_fd_sc_hd__clkbuf_2
X_2682_ _2681_/X _2532_/A _2506_/X _3171_/Q _2017_/X vssd1 vssd1 vccd1 vccd1 _2682_/X
+ sky130_fd_sc_hd__o32a_1
X_1633_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1633_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1564_ _1568_/A vssd1 vssd1 vccd1 vccd1 _1564_/Y sky130_fd_sc_hd__inv_2
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _3234_/CLK _3234_/D vssd1 vssd1 vccd1 vccd1 _3234_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3165_ _3168_/CLK _3165_/D vssd1 vssd1 vccd1 vccd1 _3165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2116_ _2905_/A _2116_/B vssd1 vssd1 vccd1 vccd1 _2116_/Y sky130_fd_sc_hd__nor2_1
X_3096_ _3100_/CLK _3096_/D vssd1 vssd1 vccd1 vccd1 _3096_/Q sky130_fd_sc_hd__dfxtp_1
X_2047_ _1857_/A _2170_/A _1880_/X _2894_/A vssd1 vssd1 vccd1 vccd1 _2047_/X sky130_fd_sc_hd__o211a_1
XFILLER_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2949_ _2962_/A vssd1 vssd1 vccd1 vccd1 _2960_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3109_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2803_ _2146_/X _2619_/C _2619_/D _1898_/X vssd1 vssd1 vccd1 vccd1 _2803_/Y sky130_fd_sc_hd__o31ai_4
X_2734_ _2835_/C _2915_/B _2734_/C _2915_/C vssd1 vssd1 vccd1 vccd1 _2736_/A sky130_fd_sc_hd__or4_1
X_2665_ _2846_/A vssd1 vssd1 vccd1 vccd1 _2665_/X sky130_fd_sc_hd__clkbuf_2
X_1616_ _1618_/A vssd1 vssd1 vccd1 vccd1 _1616_/Y sky130_fd_sc_hd__inv_2
X_2596_ _2905_/B _2885_/A _2885_/C vssd1 vssd1 vccd1 vccd1 _2596_/Y sky130_fd_sc_hd__nor3_1
XFILLER_5_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1547_ _1549_/A vssd1 vssd1 vccd1 vccd1 _1547_/Y sky130_fd_sc_hd__inv_2
X_3217_ _3234_/CLK _3217_/D vssd1 vssd1 vccd1 vccd1 _3217_/Q sky130_fd_sc_hd__dfxtp_1
X_3148_ _3152_/CLK _3148_/D vssd1 vssd1 vccd1 vccd1 _3148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_314 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_328 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3079_ _3082_/CLK _3079_/D vssd1 vssd1 vccd1 vccd1 _3079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2450_ _3112_/Q _2446_/X _2449_/X _3111_/Q vssd1 vssd1 vccd1 vccd1 _2450_/Y sky130_fd_sc_hd__a22oi_1
X_2381_ _2443_/A vssd1 vssd1 vccd1 vccd1 _2381_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3002_ _3109_/CLK _3002_/D vssd1 vssd1 vccd1 vccd1 _3002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_431 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2717_ _2766_/A vssd1 vssd1 vccd1 vccd1 _2924_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2648_ _3249_/Q vssd1 vssd1 vccd1 vccd1 _2846_/A sky130_fd_sc_hd__clkbuf_2
X_2579_ _2577_/Y _2578_/Y _2572_/X vssd1 vssd1 vccd1 vccd1 _3139_/D sky130_fd_sc_hd__a21oi_1
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_188 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1950_ _2105_/A _2105_/B vssd1 vssd1 vccd1 vccd1 _2471_/B sky130_fd_sc_hd__or2_4
X_1881_ _2170_/A _1981_/A _1880_/X _1818_/A vssd1 vssd1 vccd1 vccd1 _2137_/A sky130_fd_sc_hd__o22a_2
X_2502_ _2687_/A vssd1 vssd1 vccd1 vccd1 _2761_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2433_ _3106_/Q _2432_/X _2422_/X _3105_/Q vssd1 vssd1 vccd1 vccd1 _2433_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2364_ _2634_/A vssd1 vssd1 vccd1 vccd1 _2432_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2295_ _2280_/X _2293_/Y _2294_/X vssd1 vssd1 vccd1 vccd1 _3056_/D sky130_fd_sc_hd__a21oi_1
XFILLER_71_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3447__73 vssd1 vssd1 vccd1 vccd1 _3447__73/HI _3447_/A sky130_fd_sc_hd__conb_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_10 _3404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3375__17 vssd1 vssd1 vccd1 vccd1 _3375__17/HI _3375_/A sky130_fd_sc_hd__conb_1
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_220 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2080_ _2667_/A _2570_/C _2962_/A vssd1 vssd1 vccd1 vccd1 _2080_/X sky130_fd_sc_hd__o21a_2
XFILLER_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2982_ _3233_/CLK _2982_/D vssd1 vssd1 vccd1 vccd1 _3412_/A sky130_fd_sc_hd__dfxtp_1
X_1933_ _1933_/A vssd1 vssd1 vccd1 vccd1 _2788_/B sky130_fd_sc_hd__clkbuf_2
X_1864_ _2996_/Q _1863_/X _1783_/X _2995_/Q vssd1 vssd1 vccd1 vccd1 _1864_/Y sky130_fd_sc_hd__a22oi_1
X_1795_ _1936_/A _1858_/A _1877_/A _1953_/B vssd1 vssd1 vccd1 vccd1 _1795_/X sky130_fd_sc_hd__or4bb_2
X_3465_ _3465_/A _1644_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
X_2416_ _2443_/A vssd1 vssd1 vccd1 vccd1 _2416_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3396_ _3396_/A _1598_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2347_ _2175_/X _2346_/Y _2335_/X vssd1 vssd1 vccd1 vccd1 _3075_/D sky130_fd_sc_hd__a21oi_1
X_2278_ _3051_/Q _2271_/X _2277_/X _3050_/Q vssd1 vssd1 vccd1 vccd1 _2278_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_72_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_194 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1580_ _1580_/A vssd1 vssd1 vccd1 vccd1 _1580_/Y sky130_fd_sc_hd__inv_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3250_/CLK input2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3248_/CLK _3181_/D vssd1 vssd1 vccd1 vccd1 _3181_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2006_/Y _2231_/B _2200_/X _2048_/X vssd1 vssd1 vccd1 vccd1 _2201_/X sky130_fd_sc_hd__a31o_1
X_2132_ _2132_/A vssd1 vssd1 vccd1 vccd1 _2132_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2063_ _2198_/A _2788_/B _2492_/B vssd1 vssd1 vccd1 vccd1 _2064_/C sky130_fd_sc_hd__or3_1
X_2965_ _2971_/A _3265_/Q vssd1 vssd1 vccd1 vccd1 _2965_/X sky130_fd_sc_hd__or2_1
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2896_ _2894_/Y _2175_/C _2813_/B _2895_/X vssd1 vssd1 vccd1 vccd1 _3235_/D sky130_fd_sc_hd__o31a_1
X_1916_ _2584_/A _2835_/A _2835_/C _1916_/D vssd1 vssd1 vccd1 vccd1 _1916_/X sky130_fd_sc_hd__or4_2
X_1847_ _1895_/A _1739_/B _1845_/X _1846_/X vssd1 vssd1 vccd1 vccd1 _2477_/C sky130_fd_sc_hd__o31ai_4
Xclkbuf_leaf_25_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3233_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1778_ _2634_/A vssd1 vssd1 vccd1 vccd1 _2871_/A sky130_fd_sc_hd__clkbuf_2
X_3448_ _3448_/A _1621_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
XFILLER_76_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3379_ _3379_/A _1578_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_25_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_234 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2750_ _2750_/A _2750_/B vssd1 vssd1 vccd1 vccd1 _2751_/A sky130_fd_sc_hd__and2_1
XFILLER_8_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1701_ _3403_/A vssd1 vssd1 vccd1 vccd1 _2538_/A sky130_fd_sc_hd__clkbuf_2
X_2681_ _2681_/A _2681_/B vssd1 vssd1 vccd1 vccd1 _2681_/X sky130_fd_sc_hd__or2_1
X_1632_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1632_/Y sky130_fd_sc_hd__inv_2
X_1563_ _1575_/A vssd1 vssd1 vccd1 vccd1 _1568_/A sky130_fd_sc_hd__buf_4
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _3233_/CLK _3233_/D vssd1 vssd1 vccd1 vccd1 _3233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _3269_/CLK _3164_/D vssd1 vssd1 vccd1 vccd1 _3164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2115_ _2198_/B _2474_/B vssd1 vssd1 vccd1 vccd1 _2116_/B sky130_fd_sc_hd__nor2_1
X_3095_ _3095_/CLK _3095_/D vssd1 vssd1 vccd1 vccd1 _3095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2046_ _2046_/A _2046_/B vssd1 vssd1 vccd1 vccd1 _2046_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2948_ _1714_/X _3259_/Q _2946_/X _2947_/X vssd1 vssd1 vccd1 vccd1 _3258_/D sky130_fd_sc_hd__o211a_1
XFILLER_22_278 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2879_ _3229_/Q _2871_/X _2874_/X _3228_/Q vssd1 vssd1 vccd1 vccd1 _2879_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_38_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_45 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2802_ _2802_/A vssd1 vssd1 vccd1 vccd1 _3202_/D sky130_fd_sc_hd__clkbuf_1
X_2733_ _1696_/X _2731_/Y _2732_/X vssd1 vssd1 vccd1 vccd1 _3185_/D sky130_fd_sc_hd__o21a_1
X_2664_ _3167_/Q _2653_/X _2656_/X _3166_/Q vssd1 vssd1 vccd1 vccd1 _2664_/Y sky130_fd_sc_hd__a22oi_1
X_2595_ _2064_/X _2594_/Y _2572_/X vssd1 vssd1 vccd1 vccd1 _3143_/D sky130_fd_sc_hd__a21oi_1
X_1615_ _1618_/A vssd1 vssd1 vccd1 vccd1 _1615_/Y sky130_fd_sc_hd__inv_2
X_1546_ _1549_/A vssd1 vssd1 vccd1 vccd1 _1546_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3216_ _3234_/CLK _3216_/D vssd1 vssd1 vccd1 vccd1 _3216_/Q sky130_fd_sc_hd__dfxtp_1
X_3147_ _3152_/CLK _3147_/D vssd1 vssd1 vccd1 vccd1 _3147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_112 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3078_ _3086_/CLK _3078_/D vssd1 vssd1 vccd1 vccd1 _3078_/Q sky130_fd_sc_hd__dfxtp_1
X_2029_ _2667_/A _2915_/A _2028_/X vssd1 vssd1 vccd1 vccd1 _2029_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2380_ _2457_/A vssd1 vssd1 vccd1 vccd1 _2443_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3001_ _3105_/CLK _3001_/D vssd1 vssd1 vccd1 vccd1 _3001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2716_ _2716_/A _2716_/B vssd1 vssd1 vccd1 vccd1 _2716_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2647_ _3161_/Q _2635_/X _2642_/X _3160_/Q vssd1 vssd1 vccd1 vccd1 _2647_/Y sky130_fd_sc_hd__a22oi_1
X_2578_ _3139_/Q _2556_/X _2559_/X _3138_/Q vssd1 vssd1 vccd1 vccd1 _2578_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_200 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_454 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_468 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_90 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _1932_/A vssd1 vssd1 vccd1 vccd1 _1880_/X sky130_fd_sc_hd__clkbuf_2
X_2501_ _2973_/A _3122_/Q _1831_/X _2500_/Y vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__o22a_1
X_2432_ _2432_/A vssd1 vssd1 vccd1 vccd1 _2432_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2363_ _2892_/B _2361_/Y _2362_/X vssd1 vssd1 vccd1 vccd1 _3081_/D sky130_fd_sc_hd__a21oi_1
X_2294_ _2294_/A vssd1 vssd1 vccd1 vccd1 _2294_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_11 _3404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3462__88 vssd1 vssd1 vccd1 vccd1 _3462__88/HI _3462_/A sky130_fd_sc_hd__conb_1
XFILLER_20_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2981_ _3248_/CLK _2981_/D vssd1 vssd1 vccd1 vccd1 _3411_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1932_ _1932_/A _2026_/B vssd1 vssd1 vccd1 vccd1 _1933_/A sky130_fd_sc_hd__nor2_1
X_1863_ _2497_/A vssd1 vssd1 vccd1 vccd1 _1863_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1794_ _1794_/A vssd1 vssd1 vccd1 vccd1 _1877_/A sky130_fd_sc_hd__clkbuf_1
X_3464_ _3464_/A _1642_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
X_2415_ _3100_/Q _2403_/X _2406_/X _3099_/Q vssd1 vssd1 vccd1 vccd1 _2415_/Y sky130_fd_sc_hd__a22oi_1
X_3395_ _3395_/A _1657_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
X_2346_ _3075_/Q _2337_/X _2341_/X _3074_/Q vssd1 vssd1 vccd1 vccd1 _2346_/Y sky130_fd_sc_hd__a22oi_1
X_2277_ _2327_/A vssd1 vssd1 vccd1 vccd1 _2277_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_2_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_438 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2205_/A _2731_/A _2500_/C vssd1 vssd1 vccd1 vccd1 _2200_/X sky130_fd_sc_hd__and3_1
X_3180_ _3244_/CLK _3180_/D vssd1 vssd1 vccd1 vccd1 _3180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2131_ _2128_/Y _2552_/B _2130_/X _1992_/X vssd1 vssd1 vccd1 vccd1 _2131_/Y sky130_fd_sc_hd__o31ai_2
X_2062_ _1739_/B _1889_/X _2061_/X vssd1 vssd1 vccd1 vccd1 _2492_/B sky130_fd_sc_hd__a21o_2
XFILLER_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2964_ _2954_/X _3265_/Q _2959_/X _2963_/X vssd1 vssd1 vccd1 vccd1 _3264_/D sky130_fd_sc_hd__o211a_1
X_3432__58 vssd1 vssd1 vccd1 vccd1 _3432__58/HI _3432_/A sky130_fd_sc_hd__conb_1
X_1915_ _2901_/A _2742_/A _2079_/B vssd1 vssd1 vccd1 vccd1 _1916_/D sky130_fd_sc_hd__or3_1
X_2895_ _3235_/Q _2542_/B _2712_/X _3234_/Q _2713_/X vssd1 vssd1 vccd1 vccd1 _2895_/X
+ sky130_fd_sc_hd__o221a_1
X_1846_ _1890_/D _1877_/A _1913_/C _1858_/A vssd1 vssd1 vccd1 vccd1 _1846_/X sky130_fd_sc_hd__or4b_1
X_1777_ _2212_/A _2280_/B vssd1 vssd1 vccd1 vccd1 _1777_/Y sky130_fd_sc_hd__nand2_1
X_3447_ _3447_/A _1623_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
X_3378_ _3378_/A _1577_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
X_2329_ _2217_/Y _2328_/Y _2322_/X vssd1 vssd1 vccd1 vccd1 _3068_/D sky130_fd_sc_hd__a21oi_1
XFILLER_45_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_327 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_346 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1700_ _2959_/A vssd1 vssd1 vccd1 vccd1 _1700_/X sky130_fd_sc_hd__clkbuf_2
X_2680_ _2888_/A _2677_/X _2679_/X vssd1 vssd1 vccd1 vccd1 _3171_/D sky130_fd_sc_hd__o21a_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1631_ _1637_/A vssd1 vssd1 vccd1 vccd1 _1636_/A sky130_fd_sc_hd__buf_4
X_1562_ _1562_/A vssd1 vssd1 vccd1 vccd1 _1562_/Y sky130_fd_sc_hd__inv_2
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_191 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3232_ _3232_/CLK _3232_/D vssd1 vssd1 vccd1 vccd1 _3232_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _3269_/CLK _3163_/D vssd1 vssd1 vccd1 vccd1 _3163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2114_ _2114_/A vssd1 vssd1 vccd1 vccd1 _3022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3094_ _3095_/CLK _3094_/D vssd1 vssd1 vccd1 vccd1 _3094_/Q sky130_fd_sc_hd__dfxtp_1
X_2045_ _2537_/B _2262_/B _2045_/C vssd1 vssd1 vccd1 vccd1 _2045_/X sky130_fd_sc_hd__or3_1
XFILLER_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2947_ _2947_/A _3258_/Q vssd1 vssd1 vccd1 vccd1 _2947_/X sky130_fd_sc_hd__or2_1
X_2878_ _2792_/Y _2877_/Y _2867_/X vssd1 vssd1 vccd1 vccd1 _3228_/D sky130_fd_sc_hd__a21oi_1
X_1829_ _1895_/A vssd1 vssd1 vccd1 vccd1 _1829_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_45 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2801_ _2907_/A _2801_/B _2801_/C vssd1 vssd1 vccd1 vccd1 _2802_/A sky130_fd_sc_hd__and3_1
XFILLER_74_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2732_ _3185_/Q _2507_/X _2625_/X _3184_/Q _2678_/X vssd1 vssd1 vccd1 vccd1 _2732_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2663_ _2467_/X _2662_/Y _2649_/X vssd1 vssd1 vccd1 vccd1 _3166_/D sky130_fd_sc_hd__a21oi_1
X_2594_ _3143_/Q _2580_/X _2586_/X _3142_/Q vssd1 vssd1 vccd1 vccd1 _2594_/Y sky130_fd_sc_hd__a22oi_1
X_1614_ _1618_/A vssd1 vssd1 vccd1 vccd1 _1614_/Y sky130_fd_sc_hd__inv_2
X_1545_ _1549_/A vssd1 vssd1 vccd1 vccd1 _1545_/Y sky130_fd_sc_hd__inv_2
X_3215_ _3234_/CLK _3215_/D vssd1 vssd1 vccd1 vccd1 _3215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3146_ _3255_/CLK _3146_/D vssd1 vssd1 vccd1 vccd1 _3146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3077_ _3080_/CLK _3077_/D vssd1 vssd1 vccd1 vccd1 _3077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2028_ _2500_/A vssd1 vssd1 vccd1 vccd1 _2028_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3468__94 vssd1 vssd1 vccd1 vccd1 _3468__94/HI _3468_/A sky130_fd_sc_hd__conb_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3396__38 vssd1 vssd1 vccd1 vccd1 _3396__38/HI _3396_/A sky130_fd_sc_hd__conb_1
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_242 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3000_ _3109_/CLK _3000_/D vssd1 vssd1 vccd1 vccd1 _3000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2715_ _2710_/Y _2471_/C _2711_/X _2714_/X vssd1 vssd1 vccd1 vccd1 _3179_/D sky130_fd_sc_hd__o31a_1
X_2646_ _2041_/X _2645_/Y _2621_/X vssd1 vssd1 vccd1 vccd1 _3160_/D sky130_fd_sc_hd__a21oi_1
X_2577_ _2848_/B _2915_/A _2532_/B _2275_/X vssd1 vssd1 vccd1 vccd1 _2577_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_67_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3129_ _3154_/CLK _3129_/D vssd1 vssd1 vccd1 vccd1 _3129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2500_ _2500_/A _2500_/B _2500_/C _2500_/D vssd1 vssd1 vccd1 vccd1 _2500_/Y sky130_fd_sc_hd__nand4_1
X_2431_ _1942_/Y _2429_/Y _2430_/X vssd1 vssd1 vccd1 vccd1 _3105_/D sky130_fd_sc_hd__a21oi_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2362_ _2362_/A vssd1 vssd1 vccd1 vccd1 _2362_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2293_ _3056_/Q _2271_/X _2277_/X _3055_/Q vssd1 vssd1 vccd1 vccd1 _2293_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_2_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3230_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2629_ _2584_/X _2628_/Y _2621_/X vssd1 vssd1 vccd1 vccd1 _3155_/D sky130_fd_sc_hd__a21oi_1
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3438__64 vssd1 vssd1 vccd1 vccd1 _3438__64/HI _3438_/A sky130_fd_sc_hd__conb_1
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2980_ _3248_/CLK _2980_/D vssd1 vssd1 vccd1 vccd1 _2980_/Q sky130_fd_sc_hd__dfxtp_1
X_1931_ _1928_/Y _1930_/Y _1907_/X vssd1 vssd1 vccd1 vccd1 _3002_/D sky130_fd_sc_hd__a21oi_1
X_1862_ _1857_/Y _2667_/A _1861_/X vssd1 vssd1 vccd1 vccd1 _1862_/Y sky130_fd_sc_hd__o21ai_2
X_1793_ _3253_/Q vssd1 vssd1 vccd1 vccd1 _1858_/A sky130_fd_sc_hd__clkbuf_1
X_3463_ _3463_/A _1641_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
X_2414_ _2018_/X _2413_/X _2394_/X vssd1 vssd1 vccd1 vccd1 _3099_/D sky130_fd_sc_hd__o21a_1
X_3380__22 vssd1 vssd1 vccd1 vccd1 _3380__22/HI _3380_/A sky130_fd_sc_hd__conb_1
X_3394_ _3394_/A _1597_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
XFILLER_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2345_ _2182_/Y _2344_/Y _2335_/X vssd1 vssd1 vccd1 vccd1 _3074_/D sky130_fd_sc_hd__a21oi_1
X_2276_ _2148_/Y _2164_/X _2274_/X _2275_/X vssd1 vssd1 vccd1 vccd1 _2276_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2130_ _2223_/A _1765_/X _1991_/B _2269_/B vssd1 vssd1 vccd1 vccd1 _2130_/X sky130_fd_sc_hd__a211o_1
X_2061_ _2085_/B _2035_/B _2061_/C _2061_/D vssd1 vssd1 vccd1 vccd1 _2061_/X sky130_fd_sc_hd__and4bb_1
XFILLER_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2963_ _2971_/A _3264_/Q vssd1 vssd1 vccd1 vccd1 _2963_/X sky130_fd_sc_hd__or2_1
XFILLER_15_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1914_ _2085_/A _2026_/B _1913_/X vssd1 vssd1 vccd1 vccd1 _2079_/B sky130_fd_sc_hd__o21ai_2
X_2894_ _2894_/A _2894_/B vssd1 vssd1 vccd1 vccd1 _2894_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1845_ _1960_/B _1953_/D vssd1 vssd1 vccd1 vccd1 _1845_/X sky130_fd_sc_hd__or2b_1
X_1776_ _2537_/C _2223_/B _1765_/X _2045_/C _2731_/A vssd1 vssd1 vccd1 vccd1 _2280_/B
+ sky130_fd_sc_hd__o311a_1
X_3446_ _3446_/A _1626_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
X_3377_ _3377_/A _1576_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
X_2328_ _3068_/Q _2324_/X _2327_/X _3067_/Q vssd1 vssd1 vccd1 vccd1 _2328_/Y sky130_fd_sc_hd__a22oi_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3154_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2259_ _2046_/B _2180_/Y _2526_/A vssd1 vssd1 vccd1 vccd1 _2259_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_72_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_498 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1630_ _1630_/A vssd1 vssd1 vccd1 vccd1 _1630_/Y sky130_fd_sc_hd__inv_2
X_1561_ _1562_/A vssd1 vssd1 vccd1 vccd1 _1561_/Y sky130_fd_sc_hd__inv_2
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3231_/CLK _3231_/D vssd1 vssd1 vccd1 vccd1 _3231_/Q sky130_fd_sc_hd__dfxtp_1
X_3162_ _3268_/CLK _3162_/D vssd1 vssd1 vccd1 vccd1 _3162_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2113_ _2113_/A _2113_/B vssd1 vssd1 vccd1 vccd1 _2114_/A sky130_fd_sc_hd__and2_1
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3093_ _3095_/CLK _3093_/D vssd1 vssd1 vccd1 vccd1 _3093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2044_ _2041_/X _2042_/Y _2043_/X vssd1 vssd1 vccd1 vccd1 _3011_/D sky130_fd_sc_hd__a21oi_1
XFILLER_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2946_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2946_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2877_ _3228_/Q _2871_/X _2874_/X _3227_/Q vssd1 vssd1 vccd1 vccd1 _2877_/Y sky130_fd_sc_hd__a22oi_1
X_1828_ _1890_/D vssd1 vssd1 vccd1 vccd1 _1895_/A sky130_fd_sc_hd__buf_2
X_1759_ _1959_/A vssd1 vssd1 vccd1 vccd1 _2537_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_77_409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3429_ _3429_/A _1555_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2800_ _3202_/Q _2766_/X _2767_/X _3201_/Q vssd1 vssd1 vccd1 vccd1 _2801_/C sky130_fd_sc_hd__o22a_1
X_2731_ _2731_/A _2731_/B vssd1 vssd1 vccd1 vccd1 _2731_/Y sky130_fd_sc_hd__nand2_1
X_2662_ _3166_/Q _2653_/X _2656_/X _3165_/Q vssd1 vssd1 vccd1 vccd1 _2662_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_67_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2593_ _2498_/X _2589_/X _2592_/X _2517_/X vssd1 vssd1 vccd1 vccd1 _3142_/D sky130_fd_sc_hd__o211a_1
X_1613_ _1637_/A vssd1 vssd1 vccd1 vccd1 _1618_/A sky130_fd_sc_hd__buf_4
X_1544_ _1669_/A vssd1 vssd1 vccd1 vccd1 _1549_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3214_ _3230_/CLK _3214_/D vssd1 vssd1 vccd1 vccd1 _3214_/Q sky130_fd_sc_hd__dfxtp_1
X_3145_ _3152_/CLK _3145_/D vssd1 vssd1 vccd1 vccd1 _3145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3076_ _3080_/CLK _3076_/D vssd1 vssd1 vccd1 vccd1 _3076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2027_ _2901_/A _2778_/B _2519_/B vssd1 vssd1 vccd1 vccd1 _2915_/A sky130_fd_sc_hd__or3_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_49 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2929_ _3416_/A _2929_/B _2929_/C vssd1 vssd1 vccd1 vccd1 _2930_/A sky130_fd_sc_hd__and3_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_3_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2714_ _3179_/Q _2671_/X _2712_/X _3178_/Q _2713_/X vssd1 vssd1 vccd1 vccd1 _2714_/X
+ sky130_fd_sc_hd__o221a_1
X_2645_ _3160_/Q _2635_/X _2642_/X _3159_/Q vssd1 vssd1 vccd1 vccd1 _2645_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_10_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2576_ _2576_/A vssd1 vssd1 vccd1 vccd1 _3138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3128_ _3185_/CLK _3128_/D vssd1 vssd1 vccd1 vccd1 _3128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3059_ _3062_/CLK _3059_/D vssd1 vssd1 vccd1 vccd1 _3059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2430_ _2443_/A vssd1 vssd1 vccd1 vccd1 _2430_/X sky130_fd_sc_hd__clkbuf_2
X_2361_ _3081_/Q _2351_/X _2354_/X _3080_/Q vssd1 vssd1 vccd1 vccd1 _2361_/Y sky130_fd_sc_hd__a22oi_1
X_2292_ _2283_/X _2291_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _3055_/D sky130_fd_sc_hd__o21a_1
XFILLER_1_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2628_ _3155_/Q _2606_/X _2611_/X _3154_/Q vssd1 vssd1 vccd1 vccd1 _2628_/Y sky130_fd_sc_hd__a22oi_1
X_2559_ _2559_/A vssd1 vssd1 vccd1 vccd1 _2559_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_46 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3453__79 vssd1 vssd1 vccd1 vccd1 _3453__79/HI _3453_/A sky130_fd_sc_hd__conb_1
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1930_ _3002_/Q _1919_/X _1929_/X _3001_/Q vssd1 vssd1 vccd1 vccd1 _1930_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1861_ _2500_/A vssd1 vssd1 vccd1 vccd1 _1861_/X sky130_fd_sc_hd__buf_2
X_1792_ _3252_/Q vssd1 vssd1 vccd1 vccd1 _1936_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3462_ _3462_/A _1640_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
X_3393_ _3393_/A _1596_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
X_2413_ _3099_/Q _2497_/A _2290_/X _3098_/Q vssd1 vssd1 vccd1 vccd1 _2413_/X sky130_fd_sc_hd__a22o_1
X_2344_ _3074_/Q _2337_/X _2341_/X _3073_/Q vssd1 vssd1 vccd1 vccd1 _2344_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2275_ _2752_/A vssd1 vssd1 vccd1 vccd1 _2275_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3103_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2060_ _2905_/A _2905_/C _2742_/C vssd1 vssd1 vccd1 vccd1 _2519_/C sky130_fd_sc_hd__or3_2
X_2962_ _2962_/A vssd1 vssd1 vccd1 vccd1 _2971_/A sky130_fd_sc_hd__clkbuf_1
X_1913_ _1953_/B _1913_/B _1913_/C _1893_/B vssd1 vssd1 vccd1 vccd1 _1913_/X sky130_fd_sc_hd__or4b_2
X_2893_ _2893_/A vssd1 vssd1 vccd1 vccd1 _3234_/D sky130_fd_sc_hd__clkbuf_1
X_1844_ _2742_/A vssd1 vssd1 vccd1 vccd1 _2756_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1775_ _2788_/A _2274_/B vssd1 vssd1 vccd1 vccd1 _2731_/A sky130_fd_sc_hd__nor2_1
X_3445_ _3445_/A _1628_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3376_/A _1574_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
X_2327_ _2327_/A vssd1 vssd1 vccd1 vccd1 _2327_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2258_ _2256_/Y _2257_/Y _2241_/X vssd1 vssd1 vccd1 vccd1 _3047_/D sky130_fd_sc_hd__a21oi_1
X_2189_ _2271_/A vssd1 vssd1 vccd1 vccd1 _2189_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3423__49 vssd1 vssd1 vccd1 vccd1 _3423__49/HI _3423_/A sky130_fd_sc_hd__conb_1
XFILLER_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1560_ _1562_/A vssd1 vssd1 vccd1 vccd1 _1560_/Y sky130_fd_sc_hd__inv_2
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3230_/CLK _3230_/D vssd1 vssd1 vccd1 vccd1 _3230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _3268_/CLK _3161_/D vssd1 vssd1 vccd1 vccd1 _3161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2112_ _3022_/Q _2296_/A _2101_/A _3021_/Q _2111_/Y vssd1 vssd1 vccd1 vccd1 _2113_/B
+ sky130_fd_sc_hd__a221o_1
X_3092_ _3092_/CLK _3092_/D vssd1 vssd1 vccd1 vccd1 _3092_/Q sky130_fd_sc_hd__dfxtp_1
X_2043_ _2155_/A vssd1 vssd1 vccd1 vccd1 _2043_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2945_ _1714_/X _3258_/Q _1700_/X _2944_/X vssd1 vssd1 vccd1 vccd1 _3257_/D sky130_fd_sc_hd__o211a_1
X_2876_ _2796_/Y _2875_/Y _2867_/X vssd1 vssd1 vccd1 vccd1 _3227_/D sky130_fd_sc_hd__a21oi_1
X_1827_ _1835_/C _2747_/B vssd1 vssd1 vccd1 vccd1 _2015_/A sky130_fd_sc_hd__nor2_1
X_1758_ _2699_/A vssd1 vssd1 vccd1 vccd1 _2212_/A sky130_fd_sc_hd__buf_2
X_1689_ _3415_/A _1687_/B _1688_/Y vssd1 vssd1 vccd1 vccd1 _2985_/D sky130_fd_sc_hd__o21a_1
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3428_ _3428_/A _1554_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
XFILLER_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2730_ _2146_/X _2546_/X _2901_/C _2729_/X vssd1 vssd1 vccd1 vccd1 _3184_/D sky130_fd_sc_hd__o31a_1
X_2661_ _2638_/X _2659_/X _2660_/X _2632_/X vssd1 vssd1 vccd1 vccd1 _3165_/D sky130_fd_sc_hd__o211a_1
X_1612_ input1/X vssd1 vssd1 vccd1 vccd1 _1637_/A sky130_fd_sc_hd__clkbuf_1
X_2592_ _3142_/Q _2660_/B vssd1 vssd1 vccd1 vccd1 _2592_/X sky130_fd_sc_hd__or2_1
X_1543_ _1543_/A vssd1 vssd1 vccd1 vccd1 _1543_/Y sky130_fd_sc_hd__inv_2
X_3213_ _3230_/CLK _3213_/D vssd1 vssd1 vccd1 vccd1 _3213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3144_ _3154_/CLK _3144_/D vssd1 vssd1 vccd1 vccd1 _3144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3075_ _3194_/CLK _3075_/D vssd1 vssd1 vccd1 vccd1 _3075_/Q sky130_fd_sc_hd__dfxtp_1
X_2026_ _2094_/B _2026_/B vssd1 vssd1 vccd1 vccd1 _2519_/B sky130_fd_sc_hd__nor2_1
XFILLER_54_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2928_ _3418_/A _2704_/B _2483_/X _3245_/Q _2722_/X vssd1 vssd1 vccd1 vccd1 _3246_/D
+ sky130_fd_sc_hd__o221a_1
X_2859_ _2874_/A vssd1 vssd1 vccd1 vccd1 _2859_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_410 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3459__85 vssd1 vssd1 vccd1 vccd1 _3459__85/HI _3459_/A sky130_fd_sc_hd__conb_1
XFILLER_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3387__29 vssd1 vssd1 vccd1 vccd1 _3387__29/HI _3387_/A sky130_fd_sc_hd__conb_1
X_2713_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2713_/X sky130_fd_sc_hd__clkbuf_2
X_2644_ _2584_/X _2643_/Y _2621_/X vssd1 vssd1 vccd1 vccd1 _3159_/D sky130_fd_sc_hd__a21oi_1
X_2575_ _2769_/A _2575_/B _2575_/C vssd1 vssd1 vccd1 vccd1 _2576_/A sky130_fd_sc_hd__and3_1
XFILLER_59_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3127_ _3149_/CLK _3127_/D vssd1 vssd1 vccd1 vccd1 _3127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3058_ _3062_/CLK _3058_/D vssd1 vssd1 vccd1 vccd1 _3058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2009_ _1997_/Y _2000_/Y _2006_/Y _2008_/X _1812_/X vssd1 vssd1 vccd1 vccd1 _2009_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_332 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_70 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2360_ _2149_/Y _2359_/Y _2349_/X vssd1 vssd1 vccd1 vccd1 _3080_/D sky130_fd_sc_hd__a21oi_1
X_2291_ _3055_/Q _2081_/X _2290_/X _3054_/Q vssd1 vssd1 vccd1 vccd1 _2291_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3270_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2627_ _2667_/A _2623_/X _2626_/X vssd1 vssd1 vccd1 vccd1 _3154_/D sky130_fd_sc_hd__o21a_1
X_2558_ _1956_/X _2557_/Y _2479_/X vssd1 vssd1 vccd1 vccd1 _3133_/D sky130_fd_sc_hd__a21oi_1
X_2489_ _3120_/Q _2483_/X _2921_/A _2488_/X _2113_/A vssd1 vssd1 vccd1 vccd1 _3121_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_75_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3429__55 vssd1 vssd1 vccd1 vccd1 _3429__55/HI _3429_/A sky130_fd_sc_hd__conb_1
XFILLER_19_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1860_ _1866_/A _1935_/A _2681_/B vssd1 vssd1 vccd1 vccd1 _2667_/A sky130_fd_sc_hd__or3_4
X_1791_ _1989_/A vssd1 vssd1 vccd1 vccd1 _2026_/B sky130_fd_sc_hd__clkbuf_2
X_3461_ _3461_/A _1639_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
X_3392_ _3392_/A _1595_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_42_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2412_ _2029_/Y _2411_/Y _2401_/X vssd1 vssd1 vccd1 vccd1 _3098_/D sky130_fd_sc_hd__a21oi_1
X_2343_ _2188_/X _2342_/Y _2335_/X vssd1 vssd1 vccd1 vccd1 _3073_/D sky130_fd_sc_hd__a21oi_1
XFILLER_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2274_ _2819_/A _2274_/B _2519_/B vssd1 vssd1 vccd1 vccd1 _2274_/X sky130_fd_sc_hd__or3_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_298 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1989_ _1989_/A vssd1 vssd1 vccd1 vccd1 _2474_/B sky130_fd_sc_hd__buf_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3371__13 vssd1 vssd1 vccd1 vccd1 _3371__13/HI _3371_/A sky130_fd_sc_hd__conb_1
XFILLER_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2961_ _2954_/X _3264_/Q _2959_/X _2960_/X vssd1 vssd1 vccd1 vccd1 _3263_/D sky130_fd_sc_hd__o211a_1
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1912_ _2152_/A vssd1 vssd1 vccd1 vccd1 _2835_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2892_ _2907_/A _2892_/B _2892_/C vssd1 vssd1 vccd1 vccd1 _2893_/A sky130_fd_sc_hd__and3_1
XFILLER_8_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1843_ _1965_/A _1843_/B vssd1 vssd1 vccd1 vccd1 _2742_/A sky130_fd_sc_hd__nor2_1
X_1774_ _1924_/B _1806_/D _1947_/C _1924_/A vssd1 vssd1 vccd1 vccd1 _2274_/B sky130_fd_sc_hd__and4bb_2
X_3444_ _3444_/A _1630_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _3375_/A _1573_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
X_2326_ _2226_/Y _2325_/Y _2322_/X vssd1 vssd1 vccd1 vccd1 _3067_/D sky130_fd_sc_hd__a21oi_1
X_2257_ _3047_/Q _2244_/X _2252_/X _3046_/Q vssd1 vssd1 vccd1 vccd1 _2257_/Y sky130_fd_sc_hd__a22oi_1
X_2188_ _2894_/B _2105_/Y _1954_/X _2048_/X vssd1 vssd1 vccd1 vccd1 _2188_/X sky130_fd_sc_hd__a31o_1
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3168_/CLK _3160_/D vssd1 vssd1 vccd1 vccd1 _3160_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ _3095_/CLK _3091_/D vssd1 vssd1 vccd1 vccd1 _3091_/Q sky130_fd_sc_hd__dfxtp_1
X_2111_ _2686_/A _2537_/C vssd1 vssd1 vccd1 vccd1 _2111_/Y sky130_fd_sc_hd__nor2_1
X_2042_ _3011_/Q _1986_/X _1994_/X _3010_/Q vssd1 vssd1 vccd1 vccd1 _2042_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2944_ _2947_/A _3257_/Q vssd1 vssd1 vccd1 vccd1 _2944_/X sky130_fd_sc_hd__or2_1
XFILLER_30_282 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2875_ _3227_/Q _2871_/X _2874_/X _3226_/Q vssd1 vssd1 vccd1 vccd1 _2875_/Y sky130_fd_sc_hd__a22oi_1
X_1826_ _1949_/B vssd1 vssd1 vccd1 vccd1 _2747_/B sky130_fd_sc_hd__clkbuf_2
X_1757_ _1897_/A vssd1 vssd1 vccd1 vccd1 _2699_/A sky130_fd_sc_hd__buf_2
X_1688_ _2942_/A _2929_/C vssd1 vssd1 vccd1 vccd1 _1688_/Y sky130_fd_sc_hd__nor2_1
X_3427_ _3427_/A _1553_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _2362_/A vssd1 vssd1 vccd1 vccd1 _2309_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2660_ _3165_/Q _2660_/B vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__or2_1
X_1611_ _1611_/A vssd1 vssd1 vccd1 vccd1 _1611_/Y sky130_fd_sc_hd__inv_2
X_2591_ _2683_/A vssd1 vssd1 vccd1 vccd1 _2660_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1542_ _1543_/A vssd1 vssd1 vccd1 vccd1 _1542_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3212_ _3230_/CLK _3212_/D vssd1 vssd1 vccd1 vccd1 _3212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3143_ _3152_/CLK _3143_/D vssd1 vssd1 vccd1 vccd1 _3143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3074_ _3194_/CLK _3074_/D vssd1 vssd1 vccd1 vccd1 _3074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2025_ _2018_/X _2021_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _3009_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2927_ _2724_/Y _2926_/Y _1679_/A vssd1 vssd1 vccd1 vccd1 _3245_/D sky130_fd_sc_hd__a21oi_1
X_2858_ _2773_/X _2856_/X _2857_/X _2843_/X vssd1 vssd1 vccd1 vccd1 _3220_/D sky130_fd_sc_hd__o211a_1
X_2789_ _2540_/X _3198_/Q _2046_/B _2788_/X vssd1 vssd1 vccd1 vccd1 _2789_/X sky130_fd_sc_hd__o22a_1
X_1809_ _1935_/A _1961_/A vssd1 vssd1 vccd1 vccd1 _1896_/A sky130_fd_sc_hd__or2_1
XFILLER_49_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2712_ _2767_/A vssd1 vssd1 vccd1 vccd1 _2712_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2643_ _3159_/Q _2635_/X _2642_/X _3158_/Q vssd1 vssd1 vccd1 vccd1 _2643_/Y sky130_fd_sc_hd__a22oi_1
X_2574_ _3138_/Q _2520_/X _2522_/X _3137_/Q vssd1 vssd1 vccd1 vccd1 _2575_/C sky130_fd_sc_hd__o22a_1
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3126_ _3168_/CLK _3126_/D vssd1 vssd1 vccd1 vccd1 _3126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3057_ _3231_/CLK _3057_/D vssd1 vssd1 vccd1 vccd1 _3057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2008_ _2500_/B _1887_/B _2007_/Y vssd1 vssd1 vccd1 vccd1 _2008_/X sky130_fd_sc_hd__a21o_1
XFILLER_63_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2290_ _2874_/A vssd1 vssd1 vccd1 vccd1 _2290_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2626_ _3154_/Q _2507_/X _2625_/X _3153_/Q _2939_/B vssd1 vssd1 vccd1 vccd1 _2626_/X
+ sky130_fd_sc_hd__o221a_1
X_2557_ _3133_/Q _2556_/X _2463_/X _3132_/Q vssd1 vssd1 vccd1 vccd1 _2557_/Y sky130_fd_sc_hd__a22oi_1
X_2488_ _3121_/Q _2511_/A vssd1 vssd1 vccd1 vccd1 _2488_/X sky130_fd_sc_hd__or2_1
XFILLER_28_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3109_ _3109_/CLK _3109_/D vssd1 vssd1 vccd1 vccd1 _3109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_406 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1790_ _1794_/A _1806_/D _1888_/C vssd1 vssd1 vccd1 vccd1 _1989_/A sky130_fd_sc_hd__nand3b_1
XFILLER_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3460_ _3460_/A _1638_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
XFILLER_6_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3391_ _3391_/A _1593_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
X_2411_ _3098_/Q _2403_/X _2406_/X _3097_/Q vssd1 vssd1 vccd1 vccd1 _2411_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2342_ _3073_/Q _2337_/X _2341_/X _3072_/Q vssd1 vssd1 vccd1 vccd1 _2342_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2273_ _2270_/Y _2272_/Y _2265_/X vssd1 vssd1 vccd1 vccd1 _3050_/D sky130_fd_sc_hd__a21oi_1
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1988_ _1985_/Y _1987_/Y _1976_/X vssd1 vssd1 vccd1 vccd1 _3006_/D sky130_fd_sc_hd__a21oi_1
X_2609_ _3149_/Q _2527_/X _2533_/X _3148_/Q _2534_/X vssd1 vssd1 vccd1 vccd1 _2609_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2960_ _2960_/A _3263_/Q vssd1 vssd1 vccd1 vccd1 _2960_/X sky130_fd_sc_hd__or2_1
X_2891_ _3234_/Q _2766_/X _2767_/X _3233_/Q vssd1 vssd1 vccd1 vccd1 _2892_/C sky130_fd_sc_hd__o22a_1
X_1911_ _2122_/B vssd1 vssd1 vccd1 vccd1 _2835_/A sky130_fd_sc_hd__clkbuf_2
X_1842_ _3252_/Q _1888_/B vssd1 vssd1 vccd1 vccd1 _1965_/A sky130_fd_sc_hd__or2_2
XFILLER_8_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1773_ _3255_/Q vssd1 vssd1 vccd1 vccd1 _1806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3443_ _3443_/A _1633_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
Xrepeater3 _3248_/Q vssd1 vssd1 vccd1 vccd1 _3403_/A sky130_fd_sc_hd__clkbuf_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3374_/A _1572_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
X_2325_ _3067_/Q _2324_/X _2314_/X _3066_/Q vssd1 vssd1 vccd1 vccd1 _2325_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2256_ _2041_/C _2255_/X _2526_/A vssd1 vssd1 vccd1 vccd1 _2256_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2187_ _1804_/X _2526_/B _1829_/X vssd1 vssd1 vccd1 vccd1 _2894_/B sky130_fd_sc_hd__a21o_1
XFILLER_65_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3086_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3090_ _3092_/CLK _3090_/D vssd1 vssd1 vccd1 vccd1 _3090_/Q sky130_fd_sc_hd__dfxtp_1
X_2110_ _2108_/X _2109_/Y _2092_/X vssd1 vssd1 vccd1 vccd1 _3021_/D sky130_fd_sc_hd__a21oi_1
X_2041_ _2280_/A _2756_/C _2041_/C vssd1 vssd1 vccd1 vccd1 _2041_/X sky130_fd_sc_hd__or3_4
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_342 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2943_ _2943_/A vssd1 vssd1 vccd1 vccd1 _3256_/D sky130_fd_sc_hd__clkbuf_1
X_2874_ _2874_/A vssd1 vssd1 vccd1 vccd1 _2874_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1825_ _1836_/A _1825_/B _1888_/C vssd1 vssd1 vccd1 vccd1 _1949_/B sky130_fd_sc_hd__or3b_2
X_1756_ _1749_/Y _1755_/Y _1672_/B vssd1 vssd1 vccd1 vccd1 _2991_/D sky130_fd_sc_hd__a21oi_1
X_1687_ _3415_/A _1687_/B vssd1 vssd1 vccd1 vccd1 _2929_/C sky130_fd_sc_hd__and2_1
X_3426_ _3426_/A _1552_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _2457_/A vssd1 vssd1 vccd1 vccd1 _2362_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2239_ _1939_/Y _2710_/B _1818_/B _2760_/A _1812_/X vssd1 vssd1 vccd1 vccd1 _2239_/X
+ sky130_fd_sc_hd__a41o_2
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1610_ _1611_/A vssd1 vssd1 vccd1 vccd1 _1610_/Y sky130_fd_sc_hd__inv_2
X_2590_ _2766_/A vssd1 vssd1 vccd1 vccd1 _2683_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1541_ _1543_/A vssd1 vssd1 vccd1 vccd1 _1541_/Y sky130_fd_sc_hd__inv_2
X_3211_ _3230_/CLK _3211_/D vssd1 vssd1 vccd1 vccd1 _3211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3142_ _3154_/CLK _3142_/D vssd1 vssd1 vccd1 vccd1 _3142_/Q sky130_fd_sc_hd__dfxtp_1
X_3073_ _3080_/CLK _3073_/D vssd1 vssd1 vccd1 vccd1 _3073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2024_ _2113_/A vssd1 vssd1 vccd1 vccd1 _2024_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2926_ _3245_/Q _2019_/X _2020_/X _3244_/Q vssd1 vssd1 vccd1 vccd1 _2926_/Y sky130_fd_sc_hd__a22oi_1
X_2857_ _3220_/Q _2924_/B vssd1 vssd1 vccd1 vccd1 _2857_/X sky130_fd_sc_hd__or2_1
X_3401__43 vssd1 vssd1 vccd1 vccd1 _3401__43/HI _3401_/A sky130_fd_sc_hd__conb_1
X_1808_ _1804_/A _1947_/C _1825_/B _1924_/B vssd1 vssd1 vccd1 vccd1 _1961_/A sky130_fd_sc_hd__and4b_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2788_ _2788_/A _2788_/B _2779_/X vssd1 vssd1 vccd1 vccd1 _2788_/X sky130_fd_sc_hd__or3b_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1739_ _2223_/A _1739_/B vssd1 vssd1 vccd1 vccd1 _1739_/Y sky130_fd_sc_hd__nor2_2
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3409_ _3409_/A _1663_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2711_ _1857_/Y _2045_/C _1889_/X _2170_/C _2280_/A vssd1 vssd1 vccd1 vccd1 _2711_/X
+ sky130_fd_sc_hd__a2111o_1
X_2642_ _2783_/A vssd1 vssd1 vccd1 vccd1 _2642_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2573_ _2570_/X _2571_/Y _2572_/X vssd1 vssd1 vccd1 vccd1 _3137_/D sky130_fd_sc_hd__a21oi_1
XFILLER_59_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3125_ _3168_/CLK _3125_/D vssd1 vssd1 vccd1 vccd1 _3125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3056_ _3194_/CLK _3056_/D vssd1 vssd1 vccd1 vccd1 _3056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2007_ _2061_/D vssd1 vssd1 vccd1 vccd1 _2007_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2909_ _2885_/A _1851_/B _2760_/Y _3239_/Q _1705_/A vssd1 vssd1 vccd1 vccd1 _2909_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_58_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3464__90 vssd1 vssd1 vccd1 vccd1 _3464__90/HI _3464_/A sky130_fd_sc_hd__conb_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3392__34 vssd1 vssd1 vccd1 vccd1 _3392__34/HI _3392_/A sky130_fd_sc_hd__conb_1
XFILLER_2_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_88 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2625_ _2625_/A vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__clkbuf_2
X_2556_ _2606_/A vssd1 vssd1 vccd1 vccd1 _2556_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2487_ _2766_/A vssd1 vssd1 vccd1 vccd1 _2511_/A sky130_fd_sc_hd__clkbuf_2
X_3108_ _3109_/CLK _3108_/D vssd1 vssd1 vccd1 vccd1 _3108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3039_ _3069_/CLK _3039_/D vssd1 vssd1 vccd1 vccd1 _3039_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_37_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3253_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_418 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2410_ _2041_/X _2409_/Y _2401_/X vssd1 vssd1 vccd1 vccd1 _3097_/D sky130_fd_sc_hd__a21oi_1
X_3390_ _3390_/A _1592_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
X_2341_ _2406_/A vssd1 vssd1 vccd1 vccd1 _2341_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2272_ _3050_/Q _2271_/X _2252_/X _3049_/Q vssd1 vssd1 vccd1 vccd1 _2272_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1987_ _3006_/Q _1986_/X _1929_/X _3005_/Q vssd1 vssd1 vccd1 vccd1 _1987_/Y sky130_fd_sc_hd__a22oi_1
X_2608_ _2467_/X _2607_/Y _2600_/X vssd1 vssd1 vccd1 vccd1 _3148_/D sky130_fd_sc_hd__a21oi_1
X_2539_ _2583_/A _1939_/Y _2537_/X _2728_/B _2941_/S vssd1 vssd1 vccd1 vccd1 _2539_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_75_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3434__60 vssd1 vssd1 vccd1 vccd1 _3434__60/HI _3434_/A sky130_fd_sc_hd__conb_1
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2890_ _2212_/A _2888_/Y _2716_/Y _2889_/Y _1681_/A vssd1 vssd1 vccd1 vccd1 _3233_/D
+ sky130_fd_sc_hd__a311oi_1
X_1910_ _1910_/A vssd1 vssd1 vccd1 vccd1 _2122_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1841_ _1839_/Y _1840_/Y _1672_/B vssd1 vssd1 vccd1 vccd1 _2994_/D sky130_fd_sc_hd__a21oi_1
XFILLER_8_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1772_ _1834_/A _1959_/A _2085_/A vssd1 vssd1 vccd1 vccd1 _2788_/A sky130_fd_sc_hd__and3b_1
X_3442_ _3442_/A _1651_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
Xrepeater4 _2980_/Q vssd1 vssd1 vccd1 vccd1 _3410_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _3373_/A _1571_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2351_/A vssd1 vssd1 vccd1 vccd1 _2324_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2255_ _2170_/A _2012_/A _2036_/A _2170_/D vssd1 vssd1 vccd1 vccd1 _2255_/X sky130_fd_sc_hd__a211o_2
X_2186_ _2182_/Y _2183_/Y _2185_/X vssd1 vssd1 vccd1 vccd1 _3034_/D sky130_fd_sc_hd__a21oi_1
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_447 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_104 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2040_ _2547_/C _2693_/C _2716_/A vssd1 vssd1 vccd1 vccd1 _2041_/C sky130_fd_sc_hd__or3_2
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2942_ _2942_/A _2942_/B vssd1 vssd1 vccd1 vccd1 _2943_/A sky130_fd_sc_hd__or2_1
XFILLER_22_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_398 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2873_ _2575_/B _2872_/Y _2867_/X vssd1 vssd1 vccd1 vccd1 _3226_/D sky130_fd_sc_hd__a21oi_1
X_1824_ _1835_/C _2004_/A vssd1 vssd1 vccd1 vccd1 _2885_/A sky130_fd_sc_hd__nor2_2
X_1755_ _2991_/Q _2472_/B vssd1 vssd1 vccd1 vccd1 _1755_/Y sky130_fd_sc_hd__nand2_1
X_3364__6 vssd1 vssd1 vccd1 vccd1 _3364__6/HI _3364_/A sky130_fd_sc_hd__conb_1
X_1686_ _3414_/A _1681_/B _1685_/Y vssd1 vssd1 vccd1 vccd1 _2984_/D sky130_fd_sc_hd__o21a_1
X_3425_ _3425_/A _1549_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _3061_/Q _2297_/X _2300_/X _3060_/Q vssd1 vssd1 vccd1 vccd1 _2307_/Y sky130_fd_sc_hd__a22oi_1
X_2238_ _1739_/B _1889_/X _2061_/X vssd1 vssd1 vccd1 vccd1 _2760_/A sky130_fd_sc_hd__a21oi_1
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ _2166_/Y _2168_/Y _2155_/X vssd1 vssd1 vccd1 vccd1 _3031_/D sky130_fd_sc_hd__a21oi_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1540_ _1543_/A vssd1 vssd1 vccd1 vccd1 _1540_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3210_ _3234_/CLK _3210_/D vssd1 vssd1 vccd1 vccd1 _3210_/Q sky130_fd_sc_hd__dfxtp_1
X_3141_ _3152_/CLK _3141_/D vssd1 vssd1 vccd1 vccd1 _3141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3072_ _3080_/CLK _3072_/D vssd1 vssd1 vccd1 vccd1 _3072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2023_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2113_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2925_ _2472_/B _2923_/X _2924_/X _2722_/X vssd1 vssd1 vccd1 vccd1 _3244_/D sky130_fd_sc_hd__o211a_1
X_3398__40 vssd1 vssd1 vccd1 vccd1 _3398__40/HI _3398_/A sky130_fd_sc_hd__conb_1
X_2856_ _2905_/D _2912_/D _2164_/X _3219_/Q _1705_/A vssd1 vssd1 vccd1 vccd1 _2856_/X
+ sky130_fd_sc_hd__o32a_1
X_1807_ _1807_/A vssd1 vssd1 vccd1 vccd1 _1935_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2787_ _2217_/Y _2786_/Y _2665_/X vssd1 vssd1 vccd1 vccd1 _3198_/D sky130_fd_sc_hd__a21oi_1
X_1738_ _2267_/A vssd1 vssd1 vccd1 vccd1 _1739_/B sky130_fd_sc_hd__buf_2
X_1669_ _1669_/A vssd1 vssd1 vccd1 vccd1 _1669_/Y sky130_fd_sc_hd__inv_2
X_3408_ _3408_/A _1662_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2710_ _2710_/A _2710_/B vssd1 vssd1 vccd1 vccd1 _2710_/Y sky130_fd_sc_hd__nor2_1
X_2641_ _2638_/X _2639_/X _2640_/X _2632_/X vssd1 vssd1 vccd1 vccd1 _3158_/D sky130_fd_sc_hd__o211a_1
X_2572_ _2621_/A vssd1 vssd1 vccd1 vccd1 _2572_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3124_ _3149_/CLK _3124_/D vssd1 vssd1 vccd1 vccd1 _3124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3055_ _3194_/CLK _3055_/D vssd1 vssd1 vccd1 vccd1 _3055_/Q sky130_fd_sc_hd__dfxtp_1
X_2006_ _2710_/A _2780_/A _2005_/Y vssd1 vssd1 vccd1 vccd1 _2006_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2908_ _2908_/A vssd1 vssd1 vccd1 vccd1 _3239_/D sky130_fd_sc_hd__clkbuf_1
X_2839_ _3214_/Q _2829_/X _2832_/X _3213_/Q vssd1 vssd1 vccd1 vccd1 _2839_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3095_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3368__10 vssd1 vssd1 vccd1 vccd1 _3368__10/HI _3368_/A sky130_fd_sc_hd__conb_1
X_2624_ _2624_/A vssd1 vssd1 vccd1 vccd1 _2625_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2555_ _2555_/A vssd1 vssd1 vccd1 vccd1 _3132_/D sky130_fd_sc_hd__clkbuf_1
X_2486_ _2687_/A vssd1 vssd1 vccd1 vccd1 _2766_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3107_ _3109_/CLK _3107_/D vssd1 vssd1 vccd1 vccd1 _3107_/Q sky130_fd_sc_hd__dfxtp_1
X_3038_ _3069_/CLK _3038_/D vssd1 vssd1 vccd1 vccd1 _3038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_338 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2340_ _2585_/A vssd1 vssd1 vccd1 vccd1 _2406_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2271_ _2271_/A vssd1 vssd1 vccd1 vccd1 _2271_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1986_ _2132_/A vssd1 vssd1 vccd1 vccd1 _1986_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2607_ _3148_/Q _2606_/X _2586_/X _3147_/Q vssd1 vssd1 vccd1 vccd1 _2607_/Y sky130_fd_sc_hd__a22oi_1
X_2538_ _2538_/A vssd1 vssd1 vccd1 vccd1 _2941_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2469_ _2467_/X _2468_/Y _2458_/X vssd1 vssd1 vccd1 vccd1 _3118_/D sky130_fd_sc_hd__a21oi_1
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1840_ _2994_/Q _2773_/A _1783_/X _2993_/Q vssd1 vssd1 vccd1 vccd1 _1840_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_30_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1771_ _1953_/B vssd1 vssd1 vccd1 vccd1 _2085_/A sky130_fd_sc_hd__clkbuf_2
X_3441_ _3441_/A _1616_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
X_3372_ _3372_/A _1570_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _2232_/Y _2321_/Y _2322_/X vssd1 vssd1 vccd1 vccd1 _3066_/D sky130_fd_sc_hd__a21oi_1
XFILLER_69_146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2254_ _2249_/X _2253_/Y _2241_/X vssd1 vssd1 vccd1 vccd1 _3046_/D sky130_fd_sc_hd__a21oi_1
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2185_ _2294_/A vssd1 vssd1 vccd1 vccd1 _2185_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_388 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1969_ _2067_/A vssd1 vssd1 vccd1 vccd1 _2198_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_21_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3232_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2941_ _3256_/Q _3257_/Q _2941_/S vssd1 vssd1 vccd1 vccd1 _2942_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2872_ _3226_/Q _2871_/X _2859_/X _3225_/Q vssd1 vssd1 vccd1 vccd1 _2872_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_30_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1823_ _1823_/A vssd1 vssd1 vccd1 vccd1 _1835_/C sky130_fd_sc_hd__clkbuf_2
X_1754_ _2497_/A vssd1 vssd1 vccd1 vccd1 _2472_/B sky130_fd_sc_hd__buf_2
X_1685_ _2942_/A _1687_/B vssd1 vssd1 vccd1 vccd1 _1685_/Y sky130_fd_sc_hd__nor2_1
X_3424_ _3424_/A _1548_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _2259_/Y _2305_/Y _2294_/X vssd1 vssd1 vccd1 vccd1 _3060_/D sky130_fd_sc_hd__a21oi_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ _2235_/Y _2236_/Y _2214_/X vssd1 vssd1 vccd1 vccd1 _3043_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ _3031_/Q _2159_/X _2167_/X _3030_/Q vssd1 vssd1 vccd1 vccd1 _2168_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2099_ _2096_/X _2098_/Y _2092_/X vssd1 vssd1 vccd1 vccd1 _3019_/D sky130_fd_sc_hd__a21oi_1
XFILLER_80_174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3140_ _3152_/CLK _3140_/D vssd1 vssd1 vccd1 vccd1 _3140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3071_ _3080_/CLK _3071_/D vssd1 vssd1 vccd1 vccd1 _3071_/Q sky130_fd_sc_hd__dfxtp_1
X_2022_ _2550_/A vssd1 vssd1 vccd1 vccd1 _2713_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_399 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2924_ _3244_/Q _2924_/B vssd1 vssd1 vccd1 vccd1 _2924_/X sky130_fd_sc_hd__or2_1
X_2855_ _2810_/Y _2854_/Y _2846_/X vssd1 vssd1 vccd1 vccd1 _3219_/D sky130_fd_sc_hd__a21oi_1
X_1806_ _1888_/B _1888_/C _1836_/A _1806_/D vssd1 vssd1 vccd1 vccd1 _1807_/A sky130_fd_sc_hd__and4bb_1
X_2786_ _3198_/Q _2725_/X _2783_/X _3197_/Q vssd1 vssd1 vccd1 vccd1 _2786_/Y sky130_fd_sc_hd__a22oi_1
X_1737_ _1825_/B vssd1 vssd1 vccd1 vccd1 _2267_/A sky130_fd_sc_hd__inv_2
X_1668_ _1669_/A vssd1 vssd1 vccd1 vccd1 _1668_/Y sky130_fd_sc_hd__inv_2
X_3407_ _3407_/A _1660_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
X_1599_ _1599_/A vssd1 vssd1 vccd1 vccd1 _1599_/Y sky130_fd_sc_hd__inv_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3269_ _3269_/CLK _3269_/D vssd1 vssd1 vccd1 vccd1 _3408_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_26_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2640_ _3158_/Q _2660_/B vssd1 vssd1 vccd1 vccd1 _2640_/X sky130_fd_sc_hd__or2_1
X_2571_ _3137_/Q _2556_/X _2559_/X _3136_/Q vssd1 vssd1 vccd1 vccd1 _2571_/Y sky130_fd_sc_hd__a22oi_1
X_3123_ _3149_/CLK _3123_/D vssd1 vssd1 vccd1 vccd1 _3123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3054_ _3194_/CLK _3054_/D vssd1 vssd1 vccd1 vccd1 _3054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2005_ _2198_/B _2526_/B vssd1 vssd1 vccd1 vccd1 _2005_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2907_ _2907_/A _2907_/B _2907_/C vssd1 vssd1 vccd1 vccd1 _2908_/A sky130_fd_sc_hd__and3_1
X_2838_ _2838_/A vssd1 vssd1 vccd1 vccd1 _3213_/D sky130_fd_sc_hd__clkbuf_1
X_2769_ _2769_/A _2769_/B _2769_/C vssd1 vssd1 vccd1 vccd1 _2770_/A sky130_fd_sc_hd__and3_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3455__81 vssd1 vssd1 vccd1 vccd1 _3455__81/HI _3455_/A sky130_fd_sc_hd__conb_1
XFILLER_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2623_ _2677_/A _2623_/B _2623_/C _2623_/D vssd1 vssd1 vccd1 vccd1 _2623_/X sky130_fd_sc_hd__or4_1
X_3383__25 vssd1 vssd1 vccd1 vccd1 _3383__25/HI _3383_/A sky130_fd_sc_hd__conb_1
X_2554_ _2769_/A _2554_/B _2554_/C vssd1 vssd1 vccd1 vccd1 _2555_/A sky130_fd_sc_hd__and3_1
X_2485_ _3248_/Q _3404_/A vssd1 vssd1 vccd1 vccd1 _2687_/A sky130_fd_sc_hd__or2_1
XFILLER_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3106_ _3109_/CLK _3106_/D vssd1 vssd1 vccd1 vccd1 _3106_/Q sky130_fd_sc_hd__dfxtp_1
X_3037_ _3069_/CLK _3037_/D vssd1 vssd1 vccd1 vccd1 _3037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2270_ _2471_/C _2164_/X _2738_/D _2165_/X vssd1 vssd1 vccd1 vccd1 _2270_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_77_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1985_ _2912_/B _2912_/C _1980_/X _1984_/X _1898_/X vssd1 vssd1 vccd1 vccd1 _1985_/Y
+ sky130_fd_sc_hd__o41ai_4
X_2606_ _2606_/A vssd1 vssd1 vccd1 vccd1 _2606_/X sky130_fd_sc_hd__clkbuf_2
X_2537_ _2583_/A _2537_/B _2537_/C vssd1 vssd1 vccd1 vccd1 _2537_/X sky130_fd_sc_hd__or3_1
X_2468_ _3417_/A _2460_/X _2463_/X _3117_/Q vssd1 vssd1 vccd1 vccd1 _2468_/Y sky130_fd_sc_hd__a22oi_1
X_2399_ _2072_/Y _2398_/X _2394_/X vssd1 vssd1 vccd1 vccd1 _3093_/D sky130_fd_sc_hd__o21a_1
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_280 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3425__51 vssd1 vssd1 vccd1 vccd1 _3425__51/HI _3425_/A sky130_fd_sc_hd__conb_1
XFILLER_30_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1770_ _1823_/A vssd1 vssd1 vccd1 vccd1 _2045_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3440_ _3440_/A _1615_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
X_3371_ _3371_/A _1568_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2322_ _2362_/A vssd1 vssd1 vccd1 vccd1 _2322_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2253_ _3046_/Q _2244_/X _2252_/X _3045_/Q vssd1 vssd1 vccd1 vccd1 _2253_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_69_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2184_ _2457_/A vssd1 vssd1 vccd1 vccd1 _2294_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_334 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1968_ _1968_/A vssd1 vssd1 vccd1 vccd1 _2067_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1899_ _2157_/B _2157_/C _1898_/X vssd1 vssd1 vccd1 vccd1 _1899_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2940_ _2940_/A vssd1 vssd1 vccd1 vccd1 _3255_/D sky130_fd_sc_hd__clkbuf_1
X_2871_ _2871_/A vssd1 vssd1 vccd1 vccd1 _2871_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1822_ _2003_/A _2752_/B vssd1 vssd1 vccd1 vccd1 _2204_/A sky130_fd_sc_hd__nor2_1
X_1753_ _2634_/A vssd1 vssd1 vccd1 vccd1 _2497_/A sky130_fd_sc_hd__buf_2
X_1684_ _3413_/A _3414_/A _1684_/C vssd1 vssd1 vccd1 vccd1 _1687_/B sky130_fd_sc_hd__and3_1
X_3423_ _3423_/A _1547_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _3060_/Q _2297_/X _2300_/X _3059_/Q vssd1 vssd1 vccd1 vccd1 _2305_/Y sky130_fd_sc_hd__a22oi_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _3043_/Q _2218_/X _2227_/X _3042_/Q vssd1 vssd1 vccd1 vccd1 _2236_/Y sky130_fd_sc_hd__a22oi_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2167_ _2227_/A vssd1 vssd1 vccd1 vccd1 _2167_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_194 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2098_ _3019_/Q _2097_/X _2055_/X _3018_/Q vssd1 vssd1 vccd1 vccd1 _2098_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_80_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3070_ _3070_/CLK _3070_/D vssd1 vssd1 vccd1 vccd1 _3070_/Q sky130_fd_sc_hd__dfxtp_1
X_2021_ _3009_/Q _2019_/X _2020_/X _3008_/Q vssd1 vssd1 vccd1 vccd1 _2021_/X sky130_fd_sc_hd__a22o_1
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2923_ _2477_/A _1819_/X _2477_/C _2477_/D _2919_/X vssd1 vssd1 vccd1 vccd1 _2923_/X
+ sky130_fd_sc_hd__o41a_1
X_2854_ _3219_/Q _2853_/X _2832_/X _3218_/Q vssd1 vssd1 vccd1 vccd1 _2854_/Y sky130_fd_sc_hd__a22oi_1
X_2785_ _2217_/Y _2784_/Y _2665_/X vssd1 vssd1 vccd1 vccd1 _3197_/D sky130_fd_sc_hd__a21oi_1
X_1805_ _1932_/A _2004_/A _1804_/X vssd1 vssd1 vccd1 vccd1 _2742_/B sky130_fd_sc_hd__o21ai_4
X_1736_ _1959_/A vssd1 vssd1 vccd1 vccd1 _2223_/A sky130_fd_sc_hd__clkinv_2
X_1667_ _1669_/A vssd1 vssd1 vccd1 vccd1 _1667_/Y sky130_fd_sc_hd__inv_2
X_1598_ _1599_/A vssd1 vssd1 vccd1 vccd1 _1598_/Y sky130_fd_sc_hd__inv_2
X_3406_ _3406_/A _1659_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _3268_/CLK _3268_/D vssd1 vssd1 vccd1 vccd1 _3268_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _3040_/Q _2218_/X _2195_/X _3039_/Q vssd1 vssd1 vccd1 vccd1 _2219_/Y sky130_fd_sc_hd__a22oi_1
X_3199_ _3233_/CLK _3199_/D vssd1 vssd1 vccd1 vccd1 _3199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3389__31 vssd1 vssd1 vccd1 vccd1 _3389__31/HI _3389_/A sky130_fd_sc_hd__conb_1
XFILLER_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2570_ _2848_/A _2835_/C _2570_/C _2738_/C vssd1 vssd1 vccd1 vccd1 _2570_/X sky130_fd_sc_hd__or4_4
X_3122_ _3149_/CLK _3122_/D vssd1 vssd1 vccd1 vccd1 _3122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3053_ _3194_/CLK _3053_/D vssd1 vssd1 vccd1 vccd1 _3053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2004_ _2004_/A vssd1 vssd1 vccd1 vccd1 _2526_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2906_ _3239_/Q _2687_/X _2483_/A _3238_/Q vssd1 vssd1 vccd1 vccd1 _2907_/C sky130_fd_sc_hd__o22a_1
XFILLER_50_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2837_ _2907_/A _2837_/B _2837_/C vssd1 vssd1 vccd1 vccd1 _2838_/A sky130_fd_sc_hd__and3_1
X_2768_ _3193_/Q _2766_/X _2767_/X _3192_/Q vssd1 vssd1 vccd1 vccd1 _2769_/C sky130_fd_sc_hd__o22a_1
X_2699_ _2699_/A _3176_/Q _2699_/C vssd1 vssd1 vccd1 vccd1 _2699_/X sky130_fd_sc_hd__or3_1
X_1719_ _1794_/A vssd1 vssd1 vccd1 vccd1 _1909_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3470__96 vssd1 vssd1 vccd1 vccd1 _3470__96/HI _3470_/A sky130_fd_sc_hd__conb_1
X_2622_ _2619_/X _2620_/Y _2621_/X vssd1 vssd1 vccd1 vccd1 _3153_/D sky130_fd_sc_hd__a21oi_1
XFILLER_63_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2553_ _3132_/Q _2520_/X _2522_/X _3131_/Q vssd1 vssd1 vccd1 vccd1 _2554_/C sky130_fd_sc_hd__o22a_1
X_2484_ _2537_/C _2045_/C _1765_/X _2677_/A vssd1 vssd1 vccd1 vccd1 _2921_/A sky130_fd_sc_hd__a211o_1
X_3105_ _3105_/CLK _3105_/D vssd1 vssd1 vccd1 vccd1 _3105_/Q sky130_fd_sc_hd__dfxtp_1
X_3036_ _3080_/CLK _3036_/D vssd1 vssd1 vccd1 vccd1 _3036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3069_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_270 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1984_ _2623_/B _1997_/B _1991_/B _2552_/B vssd1 vssd1 vccd1 vccd1 _1984_/X sky130_fd_sc_hd__or4_1
XFILLER_20_159 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2605_ _2577_/Y _2604_/Y _2600_/X vssd1 vssd1 vccd1 vccd1 _3147_/D sky130_fd_sc_hd__a21oi_1
X_2536_ _2211_/B _2667_/C _2532_/X _2535_/X vssd1 vssd1 vccd1 vccd1 _3128_/D sky130_fd_sc_hd__o31a_1
X_2467_ _2467_/A _2471_/D _2885_/C vssd1 vssd1 vccd1 vccd1 _2467_/X sky130_fd_sc_hd__or3_4
XFILLER_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2398_ _3093_/Q _2081_/X _2290_/X _3092_/Q vssd1 vssd1 vccd1 vccd1 _2398_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3019_ _3092_/CLK _3019_/D vssd1 vssd1 vccd1 vccd1 _3019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_292 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3440__66 vssd1 vssd1 vccd1 vccd1 _3440__66/HI _3440_/A sky130_fd_sc_hd__conb_1
X_3370_ _3370_/A _1567_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _3066_/Q _2311_/X _2314_/X _3065_/Q vssd1 vssd1 vccd1 vccd1 _2321_/Y sky130_fd_sc_hd__a22oi_1
X_2252_ _2327_/A vssd1 vssd1 vccd1 vccd1 _2252_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2183_ _3034_/Q _2159_/X _2167_/X _3033_/Q vssd1 vssd1 vccd1 vccd1 _2183_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1967_ _2199_/B vssd1 vssd1 vccd1 vccd1 _2710_/A sky130_fd_sc_hd__clkbuf_2
X_1898_ _2752_/A vssd1 vssd1 vccd1 vccd1 _1898_/X sky130_fd_sc_hd__buf_4
X_2519_ _2738_/A _2519_/B _2519_/C _2519_/D vssd1 vssd1 vccd1 vccd1 _2524_/B sky130_fd_sc_hd__or4_1
XFILLER_68_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_88 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3268_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2870_ _2848_/X _2869_/Y _2867_/X vssd1 vssd1 vccd1 vccd1 _3225_/D sky130_fd_sc_hd__a21oi_1
X_1821_ _1843_/B vssd1 vssd1 vccd1 vccd1 _2752_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1752_ _1917_/A vssd1 vssd1 vccd1 vccd1 _2634_/A sky130_fd_sc_hd__buf_2
XFILLER_7_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1683_ _3249_/Q vssd1 vssd1 vccd1 vccd1 _2942_/A sky130_fd_sc_hd__buf_2
X_3422_ _3422_/A _1546_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _2575_/B _2303_/Y _2294_/X vssd1 vssd1 vccd1 vccd1 _3059_/D sky130_fd_sc_hd__a21oi_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _2146_/X _2072_/A _2526_/A vssd1 vssd1 vccd1 vccd1 _2235_/Y sky130_fd_sc_hd__o21ai_2
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2166_ _2742_/B _2175_/C _2164_/X _2165_/X vssd1 vssd1 vccd1 vccd1 _2166_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_53_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2097_ _2132_/A vssd1 vssd1 vccd1 vccd1 _2097_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2999_ _3105_/CLK _2999_/D vssd1 vssd1 vccd1 vccd1 _2999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_187 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2020_ _2101_/A vssd1 vssd1 vccd1 vccd1 _2020_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2922_ _2699_/C _2919_/X _2921_/Y _2843_/X vssd1 vssd1 vccd1 vccd1 _3243_/D sky130_fd_sc_hd__o211a_1
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2853_ _2871_/A vssd1 vssd1 vccd1 vccd1 _2853_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2784_ _3197_/Q _2725_/X _2783_/X _3196_/Q vssd1 vssd1 vccd1 vccd1 _2784_/Y sky130_fd_sc_hd__a22oi_1
X_1804_ _1804_/A _1947_/C _1946_/A _2058_/A vssd1 vssd1 vccd1 vccd1 _1804_/X sky130_fd_sc_hd__or4b_4
X_1735_ _1953_/D vssd1 vssd1 vccd1 vccd1 _1959_/A sky130_fd_sc_hd__clkbuf_2
X_1666_ _1666_/A vssd1 vssd1 vccd1 vccd1 _1666_/Y sky130_fd_sc_hd__inv_2
X_1597_ _1599_/A vssd1 vssd1 vccd1 vccd1 _1597_/Y sky130_fd_sc_hd__inv_2
X_3405_ _3405_/A _1658_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3267_ _3268_/CLK _3267_/D vssd1 vssd1 vccd1 vccd1 _3267_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ _2271_/A vssd1 vssd1 vccd1 vccd1 _2218_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3198_ _3233_/CLK _3198_/D vssd1 vssd1 vccd1 vccd1 _3198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2149_ _2146_/X _2532_/B _2147_/X _2148_/Y _1748_/X vssd1 vssd1 vccd1 vccd1 _2149_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3121_ _3149_/CLK _3121_/D vssd1 vssd1 vccd1 vccd1 _3121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3052_ _3070_/CLK _3052_/D vssd1 vssd1 vccd1 vccd1 _3052_/Q sky130_fd_sc_hd__dfxtp_1
X_2003_ _2003_/A vssd1 vssd1 vccd1 vccd1 _2198_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2905_ _2905_/A _2905_/B _2905_/C _2905_/D vssd1 vssd1 vccd1 vccd1 _2907_/B sky130_fd_sc_hd__or4_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2836_ _3213_/Q _2766_/X _2767_/X _3212_/Q vssd1 vssd1 vccd1 vccd1 _2837_/C sky130_fd_sc_hd__o22a_1
X_2767_ _2767_/A vssd1 vssd1 vccd1 vccd1 _2767_/X sky130_fd_sc_hd__clkbuf_2
X_1718_ _3254_/Q vssd1 vssd1 vccd1 vccd1 _1794_/A sky130_fd_sc_hd__clkbuf_1
X_2698_ _2532_/A _2848_/D _2147_/X _2915_/C _2697_/X vssd1 vssd1 vccd1 vccd1 _2698_/X
+ sky130_fd_sc_hd__o41a_1
X_1649_ _1661_/A vssd1 vssd1 vccd1 vccd1 _1654_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2621_ _2621_/A vssd1 vssd1 vccd1 vccd1 _2621_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2552_ _2681_/B _2552_/B _2552_/C _2552_/D vssd1 vssd1 vccd1 vccd1 _2554_/B sky130_fd_sc_hd__or4_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2483_ _2483_/A vssd1 vssd1 vccd1 vccd1 _2483_/X sky130_fd_sc_hd__clkbuf_2
X_3104_ _3104_/CLK _3104_/D vssd1 vssd1 vccd1 vccd1 _3104_/Q sky130_fd_sc_hd__dfxtp_1
X_3035_ _3069_/CLK _3035_/D vssd1 vssd1 vccd1 vccd1 _3035_/Q sky130_fd_sc_hd__dfxtp_1
X_3446__72 vssd1 vssd1 vccd1 vccd1 _3446__72/HI _3446_/A sky130_fd_sc_hd__conb_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2819_ _2819_/A _2819_/B _2912_/C _2819_/D vssd1 vssd1 vccd1 vccd1 _2821_/B sky130_fd_sc_hd__or4_1
XFILLER_11_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3374__16 vssd1 vssd1 vccd1 vccd1 _3374__16/HI _3374_/A sky130_fd_sc_hd__conb_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_282 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1983_ _1823_/A _1866_/A _1935_/A vssd1 vssd1 vccd1 vccd1 _2552_/B sky130_fd_sc_hd__a21o_1
X_3367__9 vssd1 vssd1 vccd1 vccd1 _3367__9/HI _3367_/A sky130_fd_sc_hd__conb_1
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2604_ _3147_/Q _2580_/X _2586_/X _3146_/Q vssd1 vssd1 vccd1 vccd1 _2604_/Y sky130_fd_sc_hd__a22oi_1
X_2535_ _3128_/Q _2527_/X _2533_/X _3127_/Q _2534_/X vssd1 vssd1 vccd1 vccd1 _2535_/X
+ sky130_fd_sc_hd__o221a_1
X_2466_ _2474_/A _2825_/A _2032_/A vssd1 vssd1 vccd1 vccd1 _2885_/C sky130_fd_sc_hd__a21o_1
X_2397_ _2076_/Y _2396_/Y _2381_/X vssd1 vssd1 vccd1 vccd1 _3092_/D sky130_fd_sc_hd__a21oi_1
XFILLER_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3018_ _3092_/CLK _3018_/D vssd1 vssd1 vccd1 vccd1 _3018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _2235_/Y _2319_/Y _2309_/X vssd1 vssd1 vccd1 vccd1 _3065_/D sky130_fd_sc_hd__a21oi_1
XFILLER_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2251_ _2585_/A vssd1 vssd1 vccd1 vccd1 _2327_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2182_ _2146_/X _2180_/Y _2619_/D _2165_/X vssd1 vssd1 vccd1 vccd1 _2182_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3116_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1966_ _2129_/B vssd1 vssd1 vccd1 vccd1 _2199_/B sky130_fd_sc_hd__clkbuf_2
X_1897_ _1897_/A vssd1 vssd1 vccd1 vccd1 _2752_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2518_ _3125_/Q _2512_/X _2516_/Y _2517_/X vssd1 vssd1 vccd1 vccd1 _3125_/D sky130_fd_sc_hd__o211a_1
X_2449_ _2559_/A vssd1 vssd1 vccd1 vccd1 _2449_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1820_ _1998_/A _1909_/A _1909_/B vssd1 vssd1 vccd1 vccd1 _1843_/B sky130_fd_sc_hd__or3_2
X_1751_ _3248_/Q _2699_/C vssd1 vssd1 vccd1 vccd1 _1917_/A sky130_fd_sc_hd__nor2_1
X_1682_ _3413_/A _1684_/C _1681_/Y vssd1 vssd1 vccd1 vccd1 _2983_/D sky130_fd_sc_hd__o21a_1
XFILLER_7_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3421_ _3421_/A _1545_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _3059_/Q _2297_/X _2300_/X _3058_/Q vssd1 vssd1 vccd1 vccd1 _2303_/Y sky130_fd_sc_hd__a22oi_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _2232_/Y _2233_/Y _2214_/X vssd1 vssd1 vccd1 vccd1 _3042_/D sky130_fd_sc_hd__a21oi_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ _2752_/A vssd1 vssd1 vccd1 vccd1 _2165_/X sky130_fd_sc_hd__buf_2
XFILLER_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2096_ _2094_/Y _2000_/Y _2731_/B _2048_/X vssd1 vssd1 vccd1 vccd1 _2096_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2998_ _3109_/CLK _2998_/D vssd1 vssd1 vccd1 vccd1 _2998_/Q sky130_fd_sc_hd__dfxtp_1
X_1949_ _1965_/A _1949_/B vssd1 vssd1 vccd1 vccd1 _2105_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_226 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2921_ _2921_/A _2921_/B vssd1 vssd1 vccd1 vccd1 _2921_/Y sky130_fd_sc_hd__nand2_1
X_2852_ _1696_/A _2180_/Y _2231_/Y _2851_/X vssd1 vssd1 vccd1 vccd1 _3218_/D sky130_fd_sc_hd__o31a_1
X_2783_ _2783_/A vssd1 vssd1 vccd1 vccd1 _2783_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1803_ _1803_/A vssd1 vssd1 vccd1 vccd1 _2004_/A sky130_fd_sc_hd__buf_2
X_1734_ _1836_/A vssd1 vssd1 vccd1 vccd1 _1953_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3404_ _3404_/A _1656_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
X_1665_ _1666_/A vssd1 vssd1 vccd1 vccd1 _1665_/Y sky130_fd_sc_hd__inv_2
X_1596_ _1599_/A vssd1 vssd1 vccd1 vccd1 _1596_/Y sky130_fd_sc_hd__inv_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3268_/CLK _3266_/D vssd1 vssd1 vccd1 vccd1 _3266_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2217_ _2477_/A _2467_/A _2471_/D _2973_/A vssd1 vssd1 vccd1 vccd1 _2217_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ _3233_/CLK _3197_/D vssd1 vssd1 vccd1 vccd1 _3197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2148_ _2128_/A _2526_/B _2566_/C vssd1 vssd1 vccd1 vccd1 _2148_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_81_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2079_ _2198_/A _2079_/B vssd1 vssd1 vccd1 vccd1 _2570_/C sky130_fd_sc_hd__or2_2
XFILLER_81_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3120_ _3154_/CLK _3120_/D vssd1 vssd1 vccd1 vccd1 _3120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3051_ _3070_/CLK _3051_/D vssd1 vssd1 vccd1 vccd1 _3051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2002_ _2825_/A vssd1 vssd1 vccd1 vccd1 _2780_/A sky130_fd_sc_hd__buf_2
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_188 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2904_ _2773_/X _2902_/X _2903_/X _2843_/X vssd1 vssd1 vccd1 vccd1 _3238_/D sky130_fd_sc_hd__o211a_1
X_2835_ _2835_/A _2905_/D _2835_/C _2566_/B vssd1 vssd1 vccd1 vccd1 _2837_/B sky130_fd_sc_hd__or4b_1
X_2766_ _2766_/A vssd1 vssd1 vccd1 vccd1 _2766_/X sky130_fd_sc_hd__clkbuf_2
X_2697_ _2941_/S _3175_/Q vssd1 vssd1 vccd1 vccd1 _2697_/X sky130_fd_sc_hd__or2_1
X_1717_ _3253_/Q vssd1 vssd1 vccd1 vccd1 _1998_/A sky130_fd_sc_hd__clkbuf_2
X_1648_ _1648_/A vssd1 vssd1 vccd1 vccd1 _1648_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _1580_/A vssd1 vssd1 vccd1 vccd1 _1579_/Y sky130_fd_sc_hd__inv_2
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3249_ _3250_/CLK hold1/X vssd1 vssd1 vccd1 vccd1 _3249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2620_ _3153_/Q _2606_/X _2611_/X _3152_/Q vssd1 vssd1 vccd1 vccd1 _2620_/Y sky130_fd_sc_hd__a22oi_1
X_2551_ _2929_/B vssd1 vssd1 vccd1 vccd1 _2769_/A sky130_fd_sc_hd__clkbuf_2
X_2482_ _2624_/A vssd1 vssd1 vccd1 vccd1 _2483_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3103_ _3103_/CLK _3103_/D vssd1 vssd1 vccd1 vccd1 _3103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3034_ _3069_/CLK _3034_/D vssd1 vssd1 vccd1 vccd1 _3034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3461__87 vssd1 vssd1 vccd1 vccd1 _3461__87/HI _3461_/A sky130_fd_sc_hd__conb_1
X_2818_ _2157_/X _2816_/Y _2817_/X vssd1 vssd1 vccd1 vccd1 _3207_/D sky130_fd_sc_hd__a21oi_1
X_2749_ _3189_/Q _2683_/A _2625_/A _3188_/Q _2393_/A vssd1 vssd1 vccd1 vccd1 _2750_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_11_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3244_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1982_ _1834_/A _1795_/X _1913_/X vssd1 vssd1 vccd1 vccd1 _1991_/B sky130_fd_sc_hd__o21ai_2
X_2603_ _2471_/B _2552_/D _2526_/Y _2602_/X vssd1 vssd1 vccd1 vccd1 _3146_/D sky130_fd_sc_hd__o31a_1
X_2534_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2534_/X sky130_fd_sc_hd__clkbuf_2
X_2465_ _1749_/Y _2464_/Y _2458_/X vssd1 vssd1 vccd1 vccd1 _3117_/D sky130_fd_sc_hd__a21oi_1
X_2396_ _3092_/Q _2383_/X _2386_/X _3091_/Q vssd1 vssd1 vccd1 vccd1 _2396_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_28_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3017_ _3092_/CLK _3017_/D vssd1 vssd1 vccd1 vccd1 _3017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _2250_/A vssd1 vssd1 vccd1 vccd1 _2585_/A sky130_fd_sc_hd__buf_2
XFILLER_77_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2181_ _2742_/B _2181_/B vssd1 vssd1 vccd1 vccd1 _2619_/D sky130_fd_sc_hd__or2_2
XFILLER_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1965_ _1965_/A vssd1 vssd1 vccd1 vccd1 _2474_/A sky130_fd_sc_hd__clkbuf_2
X_3431__57 vssd1 vssd1 vccd1 vccd1 _3431__57/HI _3431_/A sky130_fd_sc_hd__conb_1
X_1896_ _1896_/A _2152_/A _2566_/B vssd1 vssd1 vccd1 vccd1 _2157_/C sky130_fd_sc_hd__or3b_4
X_2517_ _2843_/A vssd1 vssd1 vccd1 vccd1 _2517_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2448_ _1873_/Y _2447_/Y _2443_/X vssd1 vssd1 vccd1 vccd1 _3111_/D sky130_fd_sc_hd__a21oi_1
X_2379_ _3087_/Q _2365_/X _2368_/X _3086_/Q vssd1 vssd1 vccd1 vccd1 _2379_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_24_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1750_ _3404_/A vssd1 vssd1 vccd1 vccd1 _2699_/C sky130_fd_sc_hd__clkbuf_2
X_1681_ _1681_/A _1681_/B vssd1 vssd1 vccd1 vccd1 _1681_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3420_ _3420_/A _1543_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_31_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2302_ _2270_/Y _2301_/Y _2294_/X vssd1 vssd1 vccd1 vccd1 _3058_/D sky130_fd_sc_hd__a21oi_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _3042_/Q _2218_/X _2227_/X _3041_/Q vssd1 vssd1 vccd1 vccd1 _2233_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2164_ _2738_/C vssd1 vssd1 vccd1 vccd1 _2164_/X sky130_fd_sc_hd__buf_2
X_2095_ _2223_/A _2710_/A _1831_/D _2005_/Y vssd1 vssd1 vccd1 vccd1 _2731_/B sky130_fd_sc_hd__a211oi_1
XFILLER_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2997_ _3109_/CLK _2997_/D vssd1 vssd1 vccd1 vccd1 _2997_/Q sky130_fd_sc_hd__dfxtp_1
X_1948_ _2035_/B _1947_/X _1807_/A vssd1 vssd1 vccd1 vccd1 _2105_/A sky130_fd_sc_hd__a21o_1
X_1879_ _1879_/A vssd1 vssd1 vccd1 vccd1 _2170_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2920_ _2954_/A _3242_/Q _2019_/X vssd1 vssd1 vccd1 vccd1 _2921_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2851_ _3218_/Q _2671_/X _2712_/X _3217_/Q _2713_/X vssd1 vssd1 vccd1 vccd1 _2851_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1802_ _1858_/A _1877_/A _1909_/B vssd1 vssd1 vccd1 vccd1 _1803_/A sky130_fd_sc_hd__nand3_1
X_2782_ _2778_/X _2780_/X _2781_/X vssd1 vssd1 vccd1 vccd1 _3196_/D sky130_fd_sc_hd__o21a_1
X_1733_ _3254_/Q vssd1 vssd1 vccd1 vccd1 _1836_/A sky130_fd_sc_hd__clkbuf_1
X_3403_ _3403_/A _1653_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
X_1664_ _1666_/A vssd1 vssd1 vccd1 vccd1 _1664_/Y sky130_fd_sc_hd__inv_2
X_1595_ _1599_/A vssd1 vssd1 vccd1 vccd1 _1595_/Y sky130_fd_sc_hd__inv_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3265_ _3268_/CLK _3265_/D vssd1 vssd1 vccd1 vccd1 _3265_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _2826_/A vssd1 vssd1 vccd1 vccd1 _2973_/A sky130_fd_sc_hd__buf_2
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3196_ _3241_/CLK _3196_/D vssd1 vssd1 vccd1 vccd1 _3196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2147_ _2693_/B _2693_/C _2716_/A vssd1 vssd1 vccd1 vccd1 _2147_/X sky130_fd_sc_hd__or3_2
X_2078_ _2076_/Y _2077_/Y _2043_/X vssd1 vssd1 vccd1 vccd1 _3016_/D sky130_fd_sc_hd__a21oi_1
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_14 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3467__93 vssd1 vssd1 vccd1 vccd1 _3467__93/HI _3467_/A sky130_fd_sc_hd__conb_1
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3395__37 vssd1 vssd1 vccd1 vccd1 _3395__37/HI _3395_/A sky130_fd_sc_hd__conb_1
XFILLER_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3050_ _3070_/CLK _3050_/D vssd1 vssd1 vccd1 vccd1 _3050_/Q sky130_fd_sc_hd__dfxtp_1
X_2001_ _2001_/A vssd1 vssd1 vccd1 vccd1 _2825_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2903_ _3238_/Q _2924_/B vssd1 vssd1 vccd1 vccd1 _2903_/X sky130_fd_sc_hd__or2_1
X_2834_ _2286_/X _2833_/Y _2817_/X vssd1 vssd1 vccd1 vccd1 _3212_/D sky130_fd_sc_hd__a21oi_1
X_2765_ _2765_/A _2765_/B _1939_/Y vssd1 vssd1 vccd1 vccd1 _2769_/B sky130_fd_sc_hd__or3b_1
X_1716_ _1714_/X _3408_/A _1700_/X _1715_/X vssd1 vssd1 vccd1 vccd1 _2990_/D sky130_fd_sc_hd__o211a_1
X_2696_ _2696_/A vssd1 vssd1 vccd1 vccd1 _3175_/D sky130_fd_sc_hd__clkbuf_1
X_1647_ _1648_/A vssd1 vssd1 vccd1 vccd1 _1647_/Y sky130_fd_sc_hd__inv_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _1580_/A vssd1 vssd1 vccd1 vccd1 _1578_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_215 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3248_ _3248_/CLK _3248_/D vssd1 vssd1 vccd1 vccd1 _3248_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3179_ _3241_/CLK _3179_/D vssd1 vssd1 vccd1 vccd1 _3179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_498 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2550_ _2550_/A vssd1 vssd1 vccd1 vccd1 _2929_/B sky130_fd_sc_hd__buf_2
X_2481_ _2481_/A _2699_/C vssd1 vssd1 vccd1 vccd1 _2624_/A sky130_fd_sc_hd__nand2_1
X_3102_ _3103_/CLK _3102_/D vssd1 vssd1 vccd1 vccd1 _3102_/Q sky130_fd_sc_hd__dfxtp_1
X_3033_ _3082_/CLK _3033_/D vssd1 vssd1 vccd1 vccd1 _3033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2817_ _2846_/A vssd1 vssd1 vccd1 vccd1 _2817_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2748_ _2748_/A _2813_/B _2780_/A _2075_/A vssd1 vssd1 vccd1 vccd1 _2750_/A sky130_fd_sc_hd__or4b_1
X_2679_ _3171_/Q _2507_/X _2625_/X _3170_/Q _2678_/X vssd1 vssd1 vccd1 vccd1 _2679_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3437__63 vssd1 vssd1 vccd1 vccd1 _3437__63/HI _3437_/A sky130_fd_sc_hd__conb_1
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1981_ _1981_/A _2268_/B vssd1 vssd1 vccd1 vccd1 _2623_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2602_ _3146_/Q _2527_/X _2533_/X _3145_/Q _2534_/X vssd1 vssd1 vccd1 vccd1 _2602_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2533_ _2767_/A vssd1 vssd1 vccd1 vccd1 _2533_/X sky130_fd_sc_hd__clkbuf_2
X_2464_ _3117_/Q _2460_/X _2463_/X _3116_/Q vssd1 vssd1 vccd1 vccd1 _2464_/Y sky130_fd_sc_hd__a22oi_1
X_2395_ _2080_/X _2391_/X _2394_/X vssd1 vssd1 vccd1 vccd1 _3091_/D sky130_fd_sc_hd__o21a_1
XFILLER_56_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3016_ _3092_/CLK _3016_/D vssd1 vssd1 vccd1 vccd1 _3016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_310 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2180_ _2728_/B _2180_/B vssd1 vssd1 vccd1 vccd1 _2180_/Y sky130_fd_sc_hd__nand2_2
XFILLER_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1964_ _2748_/A vssd1 vssd1 vccd1 vccd1 _2677_/B sky130_fd_sc_hd__clkbuf_2
X_1895_ _1895_/A _2012_/A vssd1 vssd1 vccd1 vccd1 _2566_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2516_ _2704_/B _2516_/B vssd1 vssd1 vccd1 vccd1 _2516_/Y sky130_fd_sc_hd__nand2_1
X_2447_ _3111_/Q _2446_/X _2435_/X _3110_/Q vssd1 vssd1 vccd1 vccd1 _2447_/Y sky130_fd_sc_hd__a22oi_1
X_2378_ _2378_/A vssd1 vssd1 vccd1 vccd1 _3086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_54 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1680_ _3413_/A _1684_/C vssd1 vssd1 vccd1 vccd1 _1681_/B sky130_fd_sc_hd__and2_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ _3058_/Q _2297_/X _2300_/X _3057_/Q vssd1 vssd1 vccd1 vccd1 _2301_/Y sky130_fd_sc_hd__a22oi_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2232_ _2888_/A _2716_/A _2231_/Y _2165_/X vssd1 vssd1 vccd1 vccd1 _2232_/Y sky130_fd_sc_hd__o31ai_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2163_ _2747_/B _2894_/A vssd1 vssd1 vccd1 vccd1 _2738_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2094_ _2677_/B _2094_/B vssd1 vssd1 vccd1 vccd1 _2094_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2996_ _3116_/CLK _2996_/D vssd1 vssd1 vccd1 vccd1 _2996_/Q sky130_fd_sc_hd__dfxtp_1
X_1947_ _1936_/A _1998_/A _1947_/C _2058_/A vssd1 vssd1 vccd1 vccd1 _1947_/X sky130_fd_sc_hd__and4bb_1
X_1878_ _1878_/A vssd1 vssd1 vccd1 vccd1 _2262_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2850_ _2848_/X _2849_/Y _2846_/X vssd1 vssd1 vccd1 vccd1 _3217_/D sky130_fd_sc_hd__a21oi_1
X_1801_ _3255_/Q vssd1 vssd1 vccd1 vccd1 _1909_/B sky130_fd_sc_hd__clkbuf_1
X_2781_ _3196_/Q _2761_/X _2625_/X _3195_/Q _2678_/X vssd1 vssd1 vccd1 vccd1 _2781_/X
+ sky130_fd_sc_hd__o221a_1
X_1732_ _1963_/A _1879_/A _1968_/A _1932_/A vssd1 vssd1 vccd1 vccd1 _2901_/A sky130_fd_sc_hd__a22o_2
X_1663_ _1666_/A vssd1 vssd1 vccd1 vccd1 _1663_/Y sky130_fd_sc_hd__inv_2
X_3402_ _3402_/A _1652_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
X_1594_ _1606_/A vssd1 vssd1 vccd1 vccd1 _1599_/A sky130_fd_sc_hd__buf_6
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _3268_/CLK _3264_/D vssd1 vssd1 vccd1 vccd1 _3264_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2215_ _2212_/Y _2213_/Y _2214_/X vssd1 vssd1 vccd1 vccd1 _3039_/D sky130_fd_sc_hd__a21oi_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _3234_/CLK _3195_/D vssd1 vssd1 vccd1 vccd1 _3195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2146_ _2756_/A vssd1 vssd1 vccd1 vccd1 _2146_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2077_ _3016_/Q _2050_/X _2055_/X _3015_/Q vssd1 vssd1 vccd1 vccd1 _2077_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2979_ _3409_/A _2212_/A _2977_/Y _2978_/X _2722_/X vssd1 vssd1 vccd1 vccd1 _3270_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3231_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_168 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2000_ _2788_/A _2778_/B vssd1 vssd1 vccd1 vccd1 _2000_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2902_ _2248_/X _2901_/Y _2699_/A _3237_/Q vssd1 vssd1 vccd1 vccd1 _2902_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2833_ _3212_/Q _2829_/X _2832_/X _3211_/Q vssd1 vssd1 vccd1 vccd1 _2833_/Y sky130_fd_sc_hd__a22oi_1
X_2764_ _1999_/A _2223_/A _1829_/X vssd1 vssd1 vccd1 vccd1 _2765_/A sky130_fd_sc_hd__a21oi_1
X_1715_ _2947_/A _3407_/A vssd1 vssd1 vccd1 vccd1 _1715_/X sky130_fd_sc_hd__or2_1
X_2695_ _2695_/A _2695_/B vssd1 vssd1 vccd1 vccd1 _2696_/A sky130_fd_sc_hd__and2_1
X_1646_ _1648_/A vssd1 vssd1 vccd1 vccd1 _1646_/Y sky130_fd_sc_hd__inv_2
X_1577_ _1580_/A vssd1 vssd1 vccd1 vccd1 _1577_/Y sky130_fd_sc_hd__inv_2
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3247_ _3248_/CLK _3247_/D vssd1 vssd1 vccd1 vccd1 _3404_/A sky130_fd_sc_hd__dfxtp_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ _3241_/CLK _3178_/D vssd1 vssd1 vccd1 vccd1 _3178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2129_ _2178_/A _2129_/B vssd1 vssd1 vccd1 vccd1 _2269_/B sky130_fd_sc_hd__nor2_1
XFILLER_54_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2480_ _2477_/X _2478_/Y _2479_/X vssd1 vssd1 vccd1 vccd1 _3120_/D sky130_fd_sc_hd__a21oi_1
X_3101_ _3104_/CLK _3101_/D vssd1 vssd1 vccd1 vccd1 _3101_/Q sky130_fd_sc_hd__dfxtp_1
X_3032_ _3082_/CLK _3032_/D vssd1 vssd1 vccd1 vccd1 _3032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2816_ _3207_/Q _2804_/X _2807_/X _3206_/Q vssd1 vssd1 vccd1 vccd1 _2816_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_11_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2747_ _3403_/A _2747_/B vssd1 vssd1 vccd1 vccd1 _2813_/B sky130_fd_sc_hd__nand2_1
X_2678_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2678_/X sky130_fd_sc_hd__clkbuf_2
X_1629_ _1630_/A vssd1 vssd1 vccd1 vccd1 _1629_/Y sky130_fd_sc_hd__inv_2
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3452__78 vssd1 vssd1 vccd1 vccd1 _3452__78/HI _3452_/A sky130_fd_sc_hd__conb_1
XFILLER_10_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3149_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_222 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1980_ _2748_/A _2105_/B _1980_/C vssd1 vssd1 vccd1 vccd1 _1980_/X sky130_fd_sc_hd__or3_1
XFILLER_41_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2601_ _2584_/X _2599_/Y _2600_/X vssd1 vssd1 vccd1 vccd1 _3145_/D sky130_fd_sc_hd__a21oi_1
XFILLER_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2532_ _2532_/A _2532_/B _2915_/C vssd1 vssd1 vccd1 vccd1 _2532_/X sky130_fd_sc_hd__or3_1
XFILLER_54_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2463_ _2559_/A vssd1 vssd1 vccd1 vccd1 _2463_/X sky130_fd_sc_hd__clkbuf_2
X_2394_ _2935_/B vssd1 vssd1 vccd1 vccd1 _2394_/X sky130_fd_sc_hd__buf_2
X_3015_ _3092_/CLK _3015_/D vssd1 vssd1 vccd1 vccd1 _3015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_447 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_99 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1963_ _1963_/A vssd1 vssd1 vccd1 vccd1 _2748_/A sky130_fd_sc_hd__clkbuf_2
X_1894_ _2004_/A _2566_/C _1940_/A vssd1 vssd1 vccd1 vccd1 _2152_/A sky130_fd_sc_hd__a21oi_2
X_2515_ _2710_/B _2248_/C _2513_/X _2514_/Y _2677_/A vssd1 vssd1 vccd1 vccd1 _2516_/B
+ sky130_fd_sc_hd__a32o_1
X_2446_ _2606_/A vssd1 vssd1 vccd1 vccd1 _2446_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2377_ _2843_/A _2377_/B vssd1 vssd1 vccd1 vccd1 _2378_/A sky130_fd_sc_hd__and2_1
XFILLER_68_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3422__48 vssd1 vssd1 vccd1 vccd1 _3422__48/HI _3422_/A sky130_fd_sc_hd__conb_1
XFILLER_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_80 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2300_ _2327_/A vssd1 vssd1 vccd1 vccd1 _2300_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2231_ _2752_/B _2231_/B vssd1 vssd1 vccd1 vccd1 _2231_/Y sky130_fd_sc_hd__nand2_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2162_ _2686_/B _2546_/C vssd1 vssd1 vccd1 vccd1 _2175_/C sky130_fd_sc_hd__or2_2
X_2093_ _2090_/Y _2091_/Y _2092_/X vssd1 vssd1 vccd1 vccd1 _3018_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2995_ _3116_/CLK _2995_/D vssd1 vssd1 vccd1 vccd1 _2995_/Q sky130_fd_sc_hd__dfxtp_1
X_1946_ _1946_/A vssd1 vssd1 vccd1 vccd1 _2035_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1877_ _1877_/A _1946_/A vssd1 vssd1 vccd1 vccd1 _1878_/A sky130_fd_sc_hd__nand2_1
X_2429_ _3105_/Q _2418_/X _2422_/X _3104_/Q vssd1 vssd1 vccd1 vccd1 _2429_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1800_ _2003_/A _2001_/A vssd1 vssd1 vccd1 vccd1 _2894_/A sky130_fd_sc_hd__nand2_2
X_2780_ _2780_/A _2885_/B _2779_/X vssd1 vssd1 vccd1 vccd1 _2780_/X sky130_fd_sc_hd__or3b_1
X_1731_ _1924_/A _2058_/A vssd1 vssd1 vccd1 vccd1 _1932_/A sky130_fd_sc_hd__or2b_2
X_1662_ _1666_/A vssd1 vssd1 vccd1 vccd1 _1662_/Y sky130_fd_sc_hd__inv_2
X_3401_ _3401_/A _1604_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
X_1593_ _1593_/A vssd1 vssd1 vccd1 vccd1 _1593_/Y sky130_fd_sc_hd__inv_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3268_/CLK _3263_/D vssd1 vssd1 vccd1 vccd1 _3263_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _2294_/A vssd1 vssd1 vccd1 vccd1 _2214_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ _3194_/CLK _3194_/D vssd1 vssd1 vccd1 vccd1 _3194_/Q sky130_fd_sc_hd__dfxtp_1
X_2145_ _2892_/B _2144_/Y _2125_/X vssd1 vssd1 vccd1 vccd1 _3027_/D sky130_fd_sc_hd__a21oi_1
XFILLER_66_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2076_ _2885_/A _1851_/B _2075_/Y _1992_/X vssd1 vssd1 vccd1 vccd1 _2076_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2978_ _2977_/A _2977_/B _2954_/A vssd1 vssd1 vccd1 vccd1 _2978_/X sky130_fd_sc_hd__a21o_1
X_1929_ _2055_/A vssd1 vssd1 vccd1 vccd1 _1929_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_386 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3458__84 vssd1 vssd1 vccd1 vccd1 _3458__84/HI _3458_/A sky130_fd_sc_hd__conb_1
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2901_ _2901_/A _2912_/B _2901_/C vssd1 vssd1 vccd1 vccd1 _2901_/Y sky130_fd_sc_hd__nor3_1
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2832_ _2874_/A vssd1 vssd1 vccd1 vccd1 _2832_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3386__28 vssd1 vssd1 vccd1 vccd1 _3386__28/HI _3386_/A sky130_fd_sc_hd__conb_1
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2763_ _1962_/X _2760_/Y _2762_/X vssd1 vssd1 vccd1 vccd1 _3192_/D sky130_fd_sc_hd__o21a_1
X_1714_ _2954_/A vssd1 vssd1 vccd1 vccd1 _1714_/X sky130_fd_sc_hd__clkbuf_2
X_2694_ _3175_/Q _2687_/X _2483_/A _3174_/Q _2508_/A vssd1 vssd1 vccd1 vccd1 _2695_/B
+ sky130_fd_sc_hd__o221a_1
X_1645_ _1648_/A vssd1 vssd1 vccd1 vccd1 _1645_/Y sky130_fd_sc_hd__inv_2
X_1576_ _1580_/A vssd1 vssd1 vccd1 vccd1 _1576_/Y sky130_fd_sc_hd__inv_2
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _3248_/CLK _3246_/D vssd1 vssd1 vccd1 vccd1 _3418_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3177_ _3233_/CLK _3177_/D vssd1 vssd1 vccd1 vccd1 _3177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2128_ _2128_/A _2710_/B vssd1 vssd1 vccd1 vccd1 _2128_/Y sky130_fd_sc_hd__nor2_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _2086_/A _1910_/A _1947_/X _2035_/B vssd1 vssd1 vccd1 vccd1 _2742_/C sky130_fd_sc_hd__a22o_1
XFILLER_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_364 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3100_ _3100_/CLK _3100_/D vssd1 vssd1 vccd1 vccd1 _3100_/Q sky130_fd_sc_hd__dfxtp_1
X_3031_ _3080_/CLK _3031_/D vssd1 vssd1 vccd1 vccd1 _3031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3255_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2815_ _2075_/Y _2819_/D _2814_/X vssd1 vssd1 vccd1 vccd1 _3206_/D sky130_fd_sc_hd__o21a_1
X_2746_ _2746_/A vssd1 vssd1 vccd1 vccd1 _3188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2677_ _2677_/A _2677_/B _2912_/B _2756_/C vssd1 vssd1 vccd1 vccd1 _2677_/X sky130_fd_sc_hd__or4_1
X_1628_ _1630_/A vssd1 vssd1 vccd1 vccd1 _1628_/Y sky130_fd_sc_hd__inv_2
X_1559_ _1562_/A vssd1 vssd1 vccd1 vccd1 _1559_/Y sky130_fd_sc_hd__inv_2
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3229_ _3230_/CLK _3229_/D vssd1 vssd1 vccd1 vccd1 _3229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3428__54 vssd1 vssd1 vccd1 vccd1 _3428__54/HI _3428_/A sky130_fd_sc_hd__conb_1
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_234 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2600_ _2621_/A vssd1 vssd1 vccd1 vccd1 _2600_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2531_ _2728_/A _2566_/B vssd1 vssd1 vccd1 vccd1 _2915_/C sky130_fd_sc_hd__nand2_1
X_2462_ _1777_/Y _2461_/Y _2458_/X vssd1 vssd1 vccd1 vccd1 _3116_/D sky130_fd_sc_hd__a21oi_1
XFILLER_47_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2393_ _2393_/A vssd1 vssd1 vccd1 vccd1 _2935_/B sky130_fd_sc_hd__clkbuf_2
X_3014_ _3095_/CLK _3014_/D vssd1 vssd1 vccd1 vccd1 _3014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2729_ _3184_/Q _2671_/X _2712_/X _3183_/Q _2713_/X vssd1 vssd1 vccd1 vccd1 _2729_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_78_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3370__12 vssd1 vssd1 vccd1 vccd1 _3370__12/HI _3370_/A sky130_fd_sc_hd__conb_1
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1962_ _2046_/A _2046_/B _2905_/A _1997_/B vssd1 vssd1 vccd1 vccd1 _1962_/X sky130_fd_sc_hd__a211o_2
X_1893_ _1913_/B _1893_/B _1913_/C _1890_/D vssd1 vssd1 vccd1 vccd1 _2566_/C sky130_fd_sc_hd__or4b_4
X_2514_ _3124_/Q vssd1 vssd1 vccd1 vccd1 _2514_/Y sky130_fd_sc_hd__inv_2
X_2445_ _2634_/A vssd1 vssd1 vccd1 vccd1 _2606_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2376_ _3086_/Q _2296_/A _2101_/A _3085_/Q _2111_/Y vssd1 vssd1 vccd1 vccd1 _2377_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_92 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2230_ _2567_/C vssd1 vssd1 vccd1 vccd1 _2888_/A sky130_fd_sc_hd__buf_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2161_ _2157_/X _2160_/Y _2155_/X vssd1 vssd1 vccd1 vccd1 _3030_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2092_ _2155_/A vssd1 vssd1 vccd1 vccd1 _2092_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2994_ _3116_/CLK _2994_/D vssd1 vssd1 vccd1 vccd1 _2994_/Q sky130_fd_sc_hd__dfxtp_1
X_1945_ _2481_/A vssd1 vssd1 vccd1 vccd1 _2738_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1876_ _1873_/Y _1875_/Y _1853_/X vssd1 vssd1 vccd1 vccd1 _2997_/D sky130_fd_sc_hd__a21oi_1
X_2428_ _1956_/X _2427_/Y _2416_/X vssd1 vssd1 vccd1 vccd1 _3104_/D sky130_fd_sc_hd__a21oi_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2359_ _3080_/Q _2351_/X _2354_/X _3079_/Q vssd1 vssd1 vccd1 vccd1 _2359_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_292 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1730_ _1888_/B vssd1 vssd1 vccd1 vccd1 _2058_/A sky130_fd_sc_hd__clkbuf_1
X_1661_ _1661_/A vssd1 vssd1 vccd1 vccd1 _1666_/A sky130_fd_sc_hd__buf_2
X_3400_ _3400_/A _1603_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
X_1592_ _1593_/A vssd1 vssd1 vccd1 vccd1 _1592_/Y sky130_fd_sc_hd__inv_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3268_/CLK _3262_/D vssd1 vssd1 vccd1 vccd1 _3262_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _3039_/Q _2189_/X _2195_/X _3038_/Q vssd1 vssd1 vccd1 vccd1 _2213_/Y sky130_fd_sc_hd__a22oi_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _3194_/CLK _3193_/D vssd1 vssd1 vccd1 vccd1 _3193_/Q sky130_fd_sc_hd__dfxtp_1
X_2144_ _3027_/Q _2132_/X _2139_/X _3026_/Q vssd1 vssd1 vccd1 vccd1 _2144_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_66_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2075_ _2075_/A _2137_/A vssd1 vssd1 vccd1 vccd1 _2075_/Y sky130_fd_sc_hd__nand2_2
XFILLER_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2977_ _2977_/A _2977_/B vssd1 vssd1 vccd1 vccd1 _2977_/Y sky130_fd_sc_hd__nor2_1
X_1928_ _1851_/B _1927_/X _1861_/X vssd1 vssd1 vccd1 vccd1 _1928_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1859_ _2085_/A _1949_/B vssd1 vssd1 vccd1 vccd1 _2681_/B sky130_fd_sc_hd__nor2_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3250_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_398 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2900_ _2041_/C _2532_/B _2885_/C _2899_/X vssd1 vssd1 vccd1 vccd1 _3237_/D sky130_fd_sc_hd__o31a_1
X_2831_ _2803_/Y _2830_/Y _2817_/X vssd1 vssd1 vccd1 vccd1 _3211_/D sky130_fd_sc_hd__a21oi_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2762_ _3192_/Q _2761_/X _2625_/X _3191_/Q _2678_/X vssd1 vssd1 vccd1 vccd1 _2762_/X
+ sky130_fd_sc_hd__o221a_1
X_1713_ _2765_/B vssd1 vssd1 vccd1 vccd1 _2954_/A sky130_fd_sc_hd__buf_2
XANTENNA_0 _2248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2693_ _2819_/A _2693_/B _2693_/C _2693_/D vssd1 vssd1 vccd1 vccd1 _2695_/A sky130_fd_sc_hd__or4_1
X_1644_ _1648_/A vssd1 vssd1 vccd1 vccd1 _1644_/Y sky130_fd_sc_hd__inv_2
X_1575_ _1575_/A vssd1 vssd1 vccd1 vccd1 _1580_/A sky130_fd_sc_hd__buf_6
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3248_/CLK _3245_/D vssd1 vssd1 vccd1 vccd1 _3245_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _3185_/CLK _3176_/D vssd1 vssd1 vccd1 vccd1 _3176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2127_ _2747_/B vssd1 vssd1 vccd1 vccd1 _2710_/B sky130_fd_sc_hd__clkbuf_2
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2058_ _2058_/A _1936_/A vssd1 vssd1 vccd1 vccd1 _2086_/A sky130_fd_sc_hd__or2b_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3030_ _3082_/CLK _3030_/D vssd1 vssd1 vccd1 vccd1 _3030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2814_ _3206_/Q _2761_/X _2528_/X _3205_/Q _2678_/X vssd1 vssd1 vccd1 vccd1 _2814_/X
+ sky130_fd_sc_hd__o221a_1
X_2745_ _2745_/A _2745_/B vssd1 vssd1 vccd1 vccd1 _2746_/A sky130_fd_sc_hd__and2_1
X_2676_ _2676_/A vssd1 vssd1 vccd1 vccd1 _3170_/D sky130_fd_sc_hd__clkbuf_1
X_1627_ _1630_/A vssd1 vssd1 vccd1 vccd1 _1627_/Y sky130_fd_sc_hd__inv_2
X_1558_ _1562_/A vssd1 vssd1 vccd1 vccd1 _1558_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3228_ _3231_/CLK _3228_/D vssd1 vssd1 vccd1 vccd1 _3228_/Q sky130_fd_sc_hd__dfxtp_1
X_3159_ _3168_/CLK _3159_/D vssd1 vssd1 vccd1 vccd1 _3159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3443__69 vssd1 vssd1 vccd1 vccd1 _3443__69/HI _3443_/A sky130_fd_sc_hd__conb_1
XFILLER_60_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2530_ _2175_/C _2742_/C _2526_/Y _2529_/X vssd1 vssd1 vccd1 vccd1 _3127_/D sky130_fd_sc_hd__o31a_1
X_2461_ _3116_/Q _2460_/X _2449_/X _3115_/Q vssd1 vssd1 vccd1 vccd1 _2461_/Y sky130_fd_sc_hd__a22oi_1
X_2392_ _2550_/A vssd1 vssd1 vccd1 vccd1 _2393_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3013_ _3013_/CLK _3013_/D vssd1 vssd1 vccd1 vccd1 _3013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2728_ _2728_/A _2728_/B vssd1 vssd1 vccd1 vccd1 _2901_/C sky130_fd_sc_hd__nand2_1
X_2659_ _2211_/B _2667_/C _2693_/D _3164_/Q _2017_/X vssd1 vssd1 vccd1 vccd1 _2659_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_47_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1961_ _1961_/A vssd1 vssd1 vccd1 vccd1 _1997_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1892_ _2756_/B _2693_/B _2038_/A vssd1 vssd1 vccd1 vccd1 _2157_/B sky130_fd_sc_hd__or3_4
X_2513_ _2474_/A _2752_/B _1897_/A _1857_/A vssd1 vssd1 vccd1 vccd1 _2513_/X sky130_fd_sc_hd__o211a_1
XFILLER_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2444_ _1882_/X _2442_/Y _2443_/X vssd1 vssd1 vccd1 vccd1 _3110_/D sky130_fd_sc_hd__a21oi_1
X_2375_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2843_/A sky130_fd_sc_hd__buf_2
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _3030_/Q _2159_/X _2139_/X _3029_/Q vssd1 vssd1 vccd1 vccd1 _2160_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2091_ _3018_/Q _2050_/X _2055_/X _3017_/Q vssd1 vssd1 vccd1 vccd1 _2091_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2993_ _3116_/CLK _2993_/D vssd1 vssd1 vccd1 vccd1 _2993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1944_ _1942_/Y _1943_/Y _1907_/X vssd1 vssd1 vccd1 vccd1 _3003_/D sky130_fd_sc_hd__a21oi_1
XFILLER_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1875_ _2997_/Q _1863_/X _1874_/X _2996_/Q vssd1 vssd1 vccd1 vccd1 _1875_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2427_ _3104_/Q _2418_/X _2422_/X _3103_/Q vssd1 vssd1 vccd1 vccd1 _2427_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2358_ _2153_/Y _2357_/Y _2349_/X vssd1 vssd1 vccd1 vccd1 _3079_/D sky130_fd_sc_hd__a21oi_1
X_2289_ _2585_/A vssd1 vssd1 vccd1 vccd1 _2874_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_411 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1660_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1660_/Y sky130_fd_sc_hd__inv_2
X_1591_ _1593_/A vssd1 vssd1 vccd1 vccd1 _1591_/Y sky130_fd_sc_hd__inv_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _3268_/CLK _3261_/D vssd1 vssd1 vccd1 vccd1 _3261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2212_ _2212_/A _2212_/B vssd1 vssd1 vccd1 vccd1 _2212_/Y sky130_fd_sc_hd__nand2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _3241_/CLK _3192_/D vssd1 vssd1 vccd1 vccd1 _3192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2143_ _2835_/A _2835_/C _2552_/C _2552_/D vssd1 vssd1 vccd1 vccd1 _2892_/B sky130_fd_sc_hd__or4_4
XFILLER_66_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2074_ _2072_/Y _2073_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _3015_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2976_ _3409_/A _3256_/Q vssd1 vssd1 vccd1 vccd1 _2977_/B sky130_fd_sc_hd__xor2_1
X_1927_ _2686_/B _2170_/C _2623_/D vssd1 vssd1 vccd1 vccd1 _1927_/X sky130_fd_sc_hd__or3_1
X_1858_ _1858_/A _1877_/A _1909_/B vssd1 vssd1 vccd1 vccd1 _1866_/A sky130_fd_sc_hd__and3_1
X_3400__42 vssd1 vssd1 vccd1 vccd1 _3400__42/HI _3400_/A sky130_fd_sc_hd__conb_1
X_1789_ _3253_/Q vssd1 vssd1 vccd1 vccd1 _1888_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3459_ _3459_/A _1636_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
XFILLER_29_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2830_ _3211_/Q _2829_/X _2807_/X _3210_/Q vssd1 vssd1 vccd1 vccd1 _2830_/Y sky130_fd_sc_hd__a22oi_1
X_2761_ _2761_/A vssd1 vssd1 vccd1 vccd1 _2761_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2692_ _2075_/Y _2181_/B _2526_/Y _2691_/X vssd1 vssd1 vccd1 vccd1 _3174_/D sky130_fd_sc_hd__o31a_1
X_1712_ _2032_/A vssd1 vssd1 vccd1 vccd1 _2765_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_1 _2575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1643_ _1661_/A vssd1 vssd1 vccd1 vccd1 _1648_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1574_ _1574_/A vssd1 vssd1 vccd1 vccd1 _1574_/Y sky130_fd_sc_hd__inv_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _3244_/CLK _3244_/D vssd1 vssd1 vccd1 vccd1 _3244_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ _3185_/CLK _3175_/D vssd1 vssd1 vccd1 vccd1 _3175_/Q sky130_fd_sc_hd__dfxtp_1
X_2126_ _2123_/Y _2124_/Y _2125_/X vssd1 vssd1 vccd1 vccd1 _3024_/D sky130_fd_sc_hd__a21oi_1
X_3449__75 vssd1 vssd1 vccd1 vccd1 _3449__75/HI _3449_/A sky130_fd_sc_hd__conb_1
XFILLER_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _2054_/Y _2056_/Y _2043_/X vssd1 vssd1 vccd1 vccd1 _3013_/D sky130_fd_sc_hd__a21oi_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3377__19 vssd1 vssd1 vccd1 vccd1 _3377__19/HI _3377_/A sky130_fd_sc_hd__conb_1
X_2959_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2959_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3391__33 vssd1 vssd1 vccd1 vccd1 _3391__33/HI _3391_/A sky130_fd_sc_hd__conb_1
XFILLER_0_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2813_ _2825_/A _2813_/B vssd1 vssd1 vccd1 vccd1 _2819_/D sky130_fd_sc_hd__or2_1
X_2744_ _3188_/Q _2683_/A _2625_/A _3187_/Q _2393_/A vssd1 vssd1 vccd1 vccd1 _2745_/B
+ sky130_fd_sc_hd__o221a_1
X_2675_ _2080_/X _2675_/B vssd1 vssd1 vccd1 vccd1 _2676_/A sky130_fd_sc_hd__and2b_1
X_1626_ _1630_/A vssd1 vssd1 vccd1 vccd1 _1626_/Y sky130_fd_sc_hd__inv_2
X_1557_ _1575_/A vssd1 vssd1 vccd1 vccd1 _1562_/A sky130_fd_sc_hd__buf_4
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3227_ _3231_/CLK _3227_/D vssd1 vssd1 vccd1 vccd1 _3227_/Q sky130_fd_sc_hd__dfxtp_1
X_3158_ _3168_/CLK _3158_/D vssd1 vssd1 vccd1 vccd1 _3158_/Q sky130_fd_sc_hd__dfxtp_1
X_2109_ _3021_/Q _2097_/X _2102_/X _3020_/Q vssd1 vssd1 vccd1 vccd1 _2109_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3089_ _3092_/CLK _3089_/D vssd1 vssd1 vccd1 vccd1 _3089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3082_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2460_ _2606_/A vssd1 vssd1 vccd1 vccd1 _2460_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2391_ _3091_/Q _2081_/X _2290_/X _3090_/Q vssd1 vssd1 vccd1 vccd1 _2391_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_200 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3012_ _3013_/CLK _3012_/D vssd1 vssd1 vccd1 vccd1 _3012_/Q sky130_fd_sc_hd__dfxtp_1
X_3419__45 vssd1 vssd1 vccd1 vccd1 _3419__45/HI _3419_/A sky130_fd_sc_hd__conb_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2727_ _2724_/Y _2726_/Y _2665_/X vssd1 vssd1 vccd1 vccd1 _3183_/D sky130_fd_sc_hd__a21oi_1
X_2658_ _2567_/X _2657_/Y _2649_/X vssd1 vssd1 vccd1 vccd1 _3164_/D sky130_fd_sc_hd__a21oi_1
X_2589_ _2248_/X _2513_/X _2540_/X _3141_/Q vssd1 vssd1 vccd1 vccd1 _2589_/X sky130_fd_sc_hd__o2bb2a_1
X_1609_ _1611_/A vssd1 vssd1 vccd1 vccd1 _1609_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1960_ _2061_/D _1960_/B _2061_/C _1960_/D vssd1 vssd1 vccd1 vccd1 _2905_/A sky130_fd_sc_hd__and4_2
XFILLER_53_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1891_ _2267_/A _1889_/X _2013_/A vssd1 vssd1 vccd1 vccd1 _2038_/A sky130_fd_sc_hd__a21o_1
X_2512_ _2704_/B vssd1 vssd1 vccd1 vccd1 _2512_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2443_ _2443_/A vssd1 vssd1 vccd1 vccd1 _2443_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2374_ _2119_/X _2373_/Y _2362_/X vssd1 vssd1 vccd1 vccd1 _3085_/D sky130_fd_sc_hd__a21oi_1
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_188 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2090_ _2848_/B _2734_/C _2532_/B _1992_/X vssd1 vssd1 vccd1 vccd1 _2090_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2992_ _3116_/CLK _2992_/D vssd1 vssd1 vccd1 vccd1 _2992_/Q sky130_fd_sc_hd__dfxtp_1
X_1943_ _3003_/Q _1919_/X _1929_/X _3002_/Q vssd1 vssd1 vccd1 vccd1 _1943_/Y sky130_fd_sc_hd__a22oi_1
X_1874_ _2055_/A vssd1 vssd1 vccd1 vccd1 _1874_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2426_ _1972_/Y _2425_/Y _2416_/X vssd1 vssd1 vccd1 vccd1 _3103_/D sky130_fd_sc_hd__a21oi_1
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2357_ _3079_/Q _2351_/X _2354_/X _3078_/Q vssd1 vssd1 vccd1 vccd1 _2357_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2288_ _2286_/X _2287_/Y _2265_/X vssd1 vssd1 vccd1 vccd1 _3054_/D sky130_fd_sc_hd__a21oi_1
XFILLER_71_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_228 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1590_ _1593_/A vssd1 vssd1 vccd1 vccd1 _1590_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3270_/CLK _3260_/D vssd1 vssd1 vccd1 vccd1 _3260_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _2825_/A _2211_/B _2467_/A _2667_/C vssd1 vssd1 vccd1 vccd1 _2212_/B sky130_fd_sc_hd__or4_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _3234_/CLK _3191_/D vssd1 vssd1 vccd1 vccd1 _3191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2142_ _2007_/Y _2067_/A _1933_/A _1934_/Y vssd1 vssd1 vccd1 vccd1 _2552_/D sky130_fd_sc_hd__a211o_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2073_ _3015_/Q _2019_/X _2020_/X _3014_/Q vssd1 vssd1 vccd1 vccd1 _2073_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2975_ _3261_/Q _3257_/Q vssd1 vssd1 vccd1 vccd1 _2977_/A sky130_fd_sc_hd__xor2_1
X_1926_ _2268_/A _2129_/B vssd1 vssd1 vccd1 vccd1 _2623_/D sky130_fd_sc_hd__nor2_1
X_1857_ _1857_/A vssd1 vssd1 vccd1 vccd1 _1857_/Y sky130_fd_sc_hd__inv_2
X_1788_ _1818_/A vssd1 vssd1 vccd1 vccd1 _2500_/B sky130_fd_sc_hd__clkbuf_2
X_3458_ _3458_/A _1635_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XFILLER_39_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3389_ _3389_/A _1591_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
X_2409_ _3097_/Q _2403_/X _2406_/X _3096_/Q vssd1 vssd1 vccd1 vccd1 _2409_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_69_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3152_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2760_ _2760_/A _2760_/B vssd1 vssd1 vccd1 vccd1 _2760_/Y sky130_fd_sc_hd__nand2_1
X_1711_ _1696_/X _3407_/A _1700_/X _1710_/X vssd1 vssd1 vccd1 vccd1 _2989_/D sky130_fd_sc_hd__o211a_1
X_2691_ _3174_/Q _2671_/X _2533_/X _3173_/Q _2534_/X vssd1 vssd1 vccd1 vccd1 _2691_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1642_ _1642_/A vssd1 vssd1 vccd1 vccd1 _1642_/Y sky130_fd_sc_hd__inv_2
XANTENNA_2 _2819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1573_ _1574_/A vssd1 vssd1 vccd1 vccd1 _1573_/Y sky130_fd_sc_hd__inv_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3244_/CLK _3243_/D vssd1 vssd1 vccd1 vccd1 _3243_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _3185_/CLK _3174_/D vssd1 vssd1 vccd1 vccd1 _3174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2125_ _2155_/A vssd1 vssd1 vccd1 vccd1 _2125_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _3013_/Q _2050_/X _2055_/X _3012_/Q vssd1 vssd1 vccd1 vccd1 _2056_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2958_ _2954_/X _3263_/Q _2946_/X _2957_/X vssd1 vssd1 vccd1 vccd1 _3262_/D sky130_fd_sc_hd__o211a_1
X_1909_ _1909_/A _1909_/B _1804_/A vssd1 vssd1 vccd1 vccd1 _1910_/A sky130_fd_sc_hd__nor3b_1
X_2889_ _3233_/Q _2511_/A _2493_/X _3232_/Q vssd1 vssd1 vccd1 vccd1 _2889_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_404 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2812_ _2810_/Y _2811_/Y _2794_/X vssd1 vssd1 vccd1 vccd1 _3205_/D sky130_fd_sc_hd__a21oi_1
X_2743_ _2765_/B _2743_/B _2743_/C vssd1 vssd1 vccd1 vccd1 _2745_/A sky130_fd_sc_hd__or3_1
X_2674_ _3170_/Q _2683_/A _2625_/A _3169_/Q _2393_/A vssd1 vssd1 vccd1 vccd1 _2675_/B
+ sky130_fd_sc_hd__o221a_1
X_1625_ _1637_/A vssd1 vssd1 vccd1 vccd1 _1630_/A sky130_fd_sc_hd__buf_4
X_1556_ _1556_/A vssd1 vssd1 vccd1 vccd1 _1556_/Y sky130_fd_sc_hd__inv_2
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _3231_/CLK _3226_/D vssd1 vssd1 vccd1 vccd1 _3226_/Q sky130_fd_sc_hd__dfxtp_1
X_3157_ _3157_/CLK _3157_/D vssd1 vssd1 vccd1 vccd1 _3157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2108_ _2105_/Y _2106_/Y _2107_/Y _2048_/X vssd1 vssd1 vccd1 vccd1 _2108_/X sky130_fd_sc_hd__a31o_1
X_3088_ _3092_/CLK _3088_/D vssd1 vssd1 vccd1 vccd1 _3088_/Q sky130_fd_sc_hd__dfxtp_1
X_2039_ _2268_/A _1981_/A _2583_/A vssd1 vssd1 vccd1 vccd1 _2716_/A sky130_fd_sc_hd__a21oi_2
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2390_ _2090_/Y _2389_/Y _2381_/X vssd1 vssd1 vccd1 vccd1 _3090_/D sky130_fd_sc_hd__a21oi_1
XFILLER_3_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3011_ _3095_/CLK _3011_/D vssd1 vssd1 vccd1 vccd1 _3011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2726_ _3183_/Q _2725_/X _2656_/X _3182_/Q vssd1 vssd1 vccd1 vccd1 _2726_/Y sky130_fd_sc_hd__a22oi_1
X_2657_ _3164_/Q _2653_/X _2656_/X _3163_/Q vssd1 vssd1 vccd1 vccd1 _2657_/Y sky130_fd_sc_hd__a22oi_1
X_1608_ _1611_/A vssd1 vssd1 vccd1 vccd1 _1608_/Y sky130_fd_sc_hd__inv_2
X_2588_ _2584_/X _2587_/Y _2572_/X vssd1 vssd1 vccd1 vccd1 _3141_/D sky130_fd_sc_hd__a21oi_1
X_1539_ _1543_/A vssd1 vssd1 vccd1 vccd1 _1539_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3209_ _3230_/CLK _3209_/D vssd1 vssd1 vccd1 vccd1 _3209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1890_ _1858_/A _1909_/B _1909_/A _1890_/D vssd1 vssd1 vccd1 vccd1 _2013_/A sky130_fd_sc_hd__and4bb_1
X_2511_ _2511_/A vssd1 vssd1 vccd1 vccd1 _2704_/B sky130_fd_sc_hd__clkbuf_2
X_2442_ _3110_/Q _2432_/X _2435_/X _3109_/Q vssd1 vssd1 vccd1 vccd1 _2442_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_45_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2373_ _3085_/Q _2365_/X _2368_/X _3084_/Q vssd1 vssd1 vccd1 vccd1 _2373_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2709_ _2638_/X _2706_/X _2707_/X _2708_/X vssd1 vssd1 vccd1 vccd1 _3178_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2991_ _3116_/CLK _2991_/D vssd1 vssd1 vccd1 vccd1 _2991_/Q sky130_fd_sc_hd__dfxtp_1
X_1942_ _2788_/B _1934_/Y _2467_/A _1941_/Y _1748_/X vssd1 vssd1 vccd1 vccd1 _1942_/Y
+ sky130_fd_sc_hd__o41ai_4
X_1873_ _2686_/C _2743_/B _1861_/X vssd1 vssd1 vccd1 vccd1 _1873_/Y sky130_fd_sc_hd__o21ai_2
X_2425_ _3103_/Q _2418_/X _2422_/X _3102_/Q vssd1 vssd1 vccd1 vccd1 _2425_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2356_ _2157_/X _2355_/Y _2349_/X vssd1 vssd1 vccd1 vccd1 _3078_/D sky130_fd_sc_hd__a21oi_1
X_2287_ _3054_/Q _2271_/X _2277_/X _3053_/Q vssd1 vssd1 vccd1 vccd1 _2287_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _1818_/A _2583_/B _1940_/A vssd1 vssd1 vccd1 vccd1 _2667_/C sky130_fd_sc_hd__a21oi_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3190_ _3244_/CLK _3190_/D vssd1 vssd1 vccd1 vccd1 _3190_/Q sky130_fd_sc_hd__dfxtp_1
X_2141_ _2138_/Y _2140_/Y _2125_/X vssd1 vssd1 vccd1 vccd1 _3026_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2072_ _2072_/A _2552_/C vssd1 vssd1 vccd1 vccd1 _2072_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2974_ _3409_/A _1696_/X _2113_/A _2973_/X vssd1 vssd1 vccd1 vccd1 _3269_/D sky130_fd_sc_hd__o211a_1
X_1925_ _1979_/B vssd1 vssd1 vccd1 vccd1 _2129_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3100_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1856_ _1856_/A vssd1 vssd1 vccd1 vccd1 _1857_/A sky130_fd_sc_hd__clkbuf_2
X_1787_ _1868_/A vssd1 vssd1 vccd1 vccd1 _1818_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3457_ _3457_/A _1634_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3388_ _3388_/A _1590_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
X_2408_ _2049_/X _2407_/Y _2401_/X vssd1 vssd1 vccd1 vccd1 _3096_/D sky130_fd_sc_hd__a21oi_1
X_2339_ _2194_/Y _2338_/Y _2335_/X vssd1 vssd1 vccd1 vccd1 _3072_/D sky130_fd_sc_hd__a21oi_1
XFILLER_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1710_ _2947_/A _3406_/A vssd1 vssd1 vccd1 vccd1 _1710_/X sky130_fd_sc_hd__or2_1
X_2690_ _2690_/A vssd1 vssd1 vccd1 vccd1 _3173_/D sky130_fd_sc_hd__clkbuf_1
X_1641_ _1642_/A vssd1 vssd1 vccd1 vccd1 _1641_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_3 _2819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1572_ _1574_/A vssd1 vssd1 vccd1 vccd1 _1572_/Y sky130_fd_sc_hd__inv_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3242_/CLK _3242_/D vssd1 vssd1 vccd1 vccd1 _3242_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _3185_/CLK _3173_/D vssd1 vssd1 vccd1 vccd1 _3173_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _3024_/Q _2097_/X _2102_/X _3023_/Q vssd1 vssd1 vccd1 vccd1 _2124_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_39_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2055_ _2055_/A vssd1 vssd1 vccd1 vccd1 _2055_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2957_ _2960_/A _3262_/Q vssd1 vssd1 vccd1 vccd1 _2957_/X sky130_fd_sc_hd__or2_1
X_1908_ _1905_/Y _1906_/Y _1907_/X vssd1 vssd1 vccd1 vccd1 _3000_/D sky130_fd_sc_hd__a21oi_1
X_2888_ _2888_/A vssd1 vssd1 vccd1 vccd1 _2888_/Y sky130_fd_sc_hd__inv_2
X_1839_ _1819_/X _1831_/X _1838_/Y _1748_/X vssd1 vssd1 vccd1 vccd1 _1839_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_77_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3454__80 vssd1 vssd1 vccd1 vccd1 _3454__80/HI _3454_/A sky130_fd_sc_hd__conb_1
X_2811_ _3205_/Q _2804_/X _2807_/X _3204_/Q vssd1 vssd1 vccd1 vccd1 _2811_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2742_ _2742_/A _2742_/B _2742_/C vssd1 vssd1 vccd1 vccd1 _2743_/C sky130_fd_sc_hd__or3_1
XFILLER_8_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2673_ _1819_/X _1851_/B _2477_/D _2672_/X vssd1 vssd1 vccd1 vccd1 _3169_/D sky130_fd_sc_hd__o31a_1
X_3382__24 vssd1 vssd1 vccd1 vccd1 _3382__24/HI _3382_/A sky130_fd_sc_hd__conb_1
X_1624_ _1624_/A vssd1 vssd1 vccd1 vccd1 _1624_/Y sky130_fd_sc_hd__inv_2
X_1555_ _1556_/A vssd1 vssd1 vccd1 vccd1 _1555_/Y sky130_fd_sc_hd__inv_2
X_3225_ _3231_/CLK _3225_/D vssd1 vssd1 vccd1 vccd1 _3225_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3156_ _3157_/CLK _3156_/D vssd1 vssd1 vccd1 vccd1 _3156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2107_ _2211_/B _2170_/C _2623_/D vssd1 vssd1 vccd1 vccd1 _2107_/Y sky130_fd_sc_hd__nor3_1
XFILLER_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3087_ _3092_/CLK _3087_/D vssd1 vssd1 vccd1 vccd1 _3087_/Q sky130_fd_sc_hd__dfxtp_1
X_2038_ _2038_/A vssd1 vssd1 vccd1 vccd1 _2693_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_42_408 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_14 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3234_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_88 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3010_ _3100_/CLK _3010_/D vssd1 vssd1 vccd1 vccd1 _3010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2725_ _2829_/A vssd1 vssd1 vccd1 vccd1 _2725_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2656_ _2783_/A vssd1 vssd1 vccd1 vccd1 _2656_/X sky130_fd_sc_hd__clkbuf_2
X_1607_ _1611_/A vssd1 vssd1 vccd1 vccd1 _1607_/Y sky130_fd_sc_hd__inv_2
X_2587_ _3141_/Q _2580_/X _2586_/X _3140_/Q vssd1 vssd1 vccd1 vccd1 _2587_/Y sky130_fd_sc_hd__a22oi_1
X_1538_ _1669_/A vssd1 vssd1 vccd1 vccd1 _1543_/A sky130_fd_sc_hd__buf_2
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3208_ _3234_/CLK _3208_/D vssd1 vssd1 vccd1 vccd1 _3208_/Q sky130_fd_sc_hd__dfxtp_1
X_3139_ _3152_/CLK _3139_/D vssd1 vssd1 vccd1 vccd1 _3139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3424__50 vssd1 vssd1 vccd1 vccd1 _3424__50/HI _3424_/A sky130_fd_sc_hd__conb_1
X_2510_ _2255_/X _2506_/X _2509_/X vssd1 vssd1 vccd1 vccd1 _3124_/D sky130_fd_sc_hd__o21a_1
X_2441_ _1899_/Y _2440_/Y _2430_/X vssd1 vssd1 vccd1 vccd1 _3109_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2372_ _2123_/Y _2371_/Y _2362_/X vssd1 vssd1 vccd1 vccd1 _3084_/D sky130_fd_sc_hd__a21oi_1
XFILLER_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2708_ _2843_/A vssd1 vssd1 vccd1 vccd1 _2708_/X sky130_fd_sc_hd__clkbuf_2
X_2639_ _2973_/A _3157_/Q _2157_/B _2693_/D vssd1 vssd1 vccd1 vccd1 _2639_/X sky130_fd_sc_hd__o22a_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_190 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2990_ _3253_/CLK _2990_/D vssd1 vssd1 vccd1 vccd1 _3407_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1941_ _1939_/Y _2752_/B _2046_/A vssd1 vssd1 vccd1 vccd1 _1941_/Y sky130_fd_sc_hd__a21oi_1
X_1872_ _2546_/C _2075_/A vssd1 vssd1 vccd1 vccd1 _2743_/B sky130_fd_sc_hd__or2b_1
X_2424_ _1985_/Y _2423_/Y _2416_/X vssd1 vssd1 vccd1 vccd1 _3102_/D sky130_fd_sc_hd__a21oi_1
X_2355_ _3078_/Q _2351_/X _2354_/X _3077_/Q vssd1 vssd1 vccd1 vccd1 _2355_/Y sky130_fd_sc_hd__a22oi_1
X_2286_ _2105_/Y _2106_/Y _1954_/X _2280_/A vssd1 vssd1 vccd1 vccd1 _2286_/X sky130_fd_sc_hd__a31o_2
XFILLER_37_396 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2140_ _3026_/Q _2132_/X _2139_/X _3025_/Q vssd1 vssd1 vccd1 vccd1 _2140_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2071_ _2198_/B _2001_/A _2032_/A vssd1 vssd1 vccd1 vccd1 _2552_/C sky130_fd_sc_hd__a21o_1
XFILLER_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2973_ _2973_/A _3408_/A vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__or2_1
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1924_ _1924_/A _1924_/B vssd1 vssd1 vccd1 vccd1 _1979_/B sky130_fd_sc_hd__and2_1
X_1855_ _1953_/D _1960_/D vssd1 vssd1 vccd1 vccd1 _1856_/A sky130_fd_sc_hd__or2b_1
X_1786_ _3253_/Q _1794_/A _1806_/D vssd1 vssd1 vccd1 vccd1 _1868_/A sky130_fd_sc_hd__or3b_1
X_3456_ _3456_/A _1632_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
X_3387_ _3387_/A _1589_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
X_2407_ _3096_/Q _2403_/X _2406_/X _3095_/Q vssd1 vssd1 vccd1 vccd1 _2407_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_57_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2338_ _3072_/Q _2337_/X _2327_/X _3071_/Q vssd1 vssd1 vccd1 vccd1 _2338_/Y sky130_fd_sc_hd__a22oi_1
X_2269_ _2819_/B _2269_/B _2912_/C _2269_/D vssd1 vssd1 vccd1 vccd1 _2738_/D sky130_fd_sc_hd__or4_2
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3388__30 vssd1 vssd1 vccd1 vccd1 _3388__30/HI _3388_/A sky130_fd_sc_hd__conb_1
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1640_ _1642_/A vssd1 vssd1 vccd1 vccd1 _1640_/Y sky130_fd_sc_hd__inv_2
X_1571_ _1574_/A vssd1 vssd1 vccd1 vccd1 _1571_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_4 _2843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3241_/CLK _3241_/D vssd1 vssd1 vccd1 vccd1 _3241_/Q sky130_fd_sc_hd__dfxtp_1
X_3172_ _3185_/CLK _3172_/D vssd1 vssd1 vccd1 vccd1 _3172_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _2623_/C _2122_/X _2028_/X vssd1 vssd1 vccd1 vccd1 _2123_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_222 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2054_ _1934_/Y _2053_/X _2028_/X vssd1 vssd1 vccd1 vccd1 _2054_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2956_ _2954_/X _3262_/Q _2946_/X _2955_/X vssd1 vssd1 vccd1 vccd1 _3261_/D sky130_fd_sc_hd__o211a_1
X_1907_ _2942_/A vssd1 vssd1 vccd1 vccd1 _1907_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2887_ _2180_/Y _2885_/X _2886_/X vssd1 vssd1 vccd1 vccd1 _3232_/D sky130_fd_sc_hd__o21a_1
X_1838_ _1838_/A _1887_/B vssd1 vssd1 vccd1 vccd1 _1838_/Y sky130_fd_sc_hd__nand2_1
X_1769_ _1951_/B vssd1 vssd1 vccd1 vccd1 _1823_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3439_ _3439_/A _1614_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_314 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_262 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2810_ _2584_/B _2693_/C _2584_/D _2017_/X vssd1 vssd1 vccd1 vccd1 _2810_/Y sky130_fd_sc_hd__o31ai_4
X_2741_ _2741_/A vssd1 vssd1 vccd1 vccd1 _3187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2672_ _3169_/Q _2671_/X _2533_/X _3168_/Q _2534_/X vssd1 vssd1 vccd1 vccd1 _2672_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1623_ _1624_/A vssd1 vssd1 vccd1 vccd1 _1623_/Y sky130_fd_sc_hd__inv_2
X_1554_ _1556_/A vssd1 vssd1 vccd1 vccd1 _1554_/Y sky130_fd_sc_hd__inv_2
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3224_ _3231_/CLK _3224_/D vssd1 vssd1 vccd1 vccd1 _3224_/Q sky130_fd_sc_hd__dfxtp_1
.ends

